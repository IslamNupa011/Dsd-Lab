CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
64
13 Logic Switch~
5 334 2102 0 1 11
0 58
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 s2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9796 0 0
2
43495 0
0
13 Logic Switch~
5 202 2111 0 10 11
0 59 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 s1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5952 0 0
2
43495 0
0
13 Logic Switch~
5 75 2116 0 1 11
0 61
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 s0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3649 0 0
2
43495 0
0
13 Logic Switch~
5 389 40 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
2 a0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3716 0 0
2
43495 0
0
13 Logic Switch~
5 282 45 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 a1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4797 0 0
2
43495 0
0
13 Logic Switch~
5 156 46 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 a2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4681 0 0
2
43495 0
0
13 Logic Switch~
5 41 50 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 a3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9730 0 0
2
43495 0
0
2 +V
167 887 584 0 1 3
0 7
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9874 0 0
2
43495.1 0
0
7 Ground~
168 884 494 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
364 0 0
2
43495.1 0
0
5 4049~
219 80 26 0 2 22
0 6 8
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U23A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 23 0
1 U
3656 0 0
2
43495 0
0
5 4049~
219 200 25 0 2 22
0 3 9
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 17 0
1 U
3131 0 0
2
43495 0
0
5 4049~
219 319 16 0 2 22
0 4 11
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 17 0
1 U
6772 0 0
2
43495 0
0
5 4049~
219 441 12 0 2 22
0 5 13
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 17 0
1 U
9557 0 0
2
43495 0
0
8 4-In OR~
219 737 1921 0 5 22
0 19 18 17 16 15
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U22B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 22 0
1 U
5789 0 0
2
43495 0
0
8 4-In OR~
219 729 1670 0 5 22
0 24 23 22 21 20
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U22A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 22 0
1 U
7328 0 0
2
43495 0
0
5 4071~
219 926 1796 0 3 22
0 20 15 14
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U19D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 19 0
1 U
4799 0 0
2
43495 0
0
5 4071~
219 892 1276 0 3 22
0 31 26 25
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U19C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 19 0
1 U
9196 0 0
2
43495 0
0
8 4-In OR~
219 745 1405 0 5 22
0 30 29 28 27 26
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U21B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 21 0
1 U
3857 0 0
2
43495 0
0
8 4-In OR~
219 742 1181 0 5 22
0 35 34 33 32 31
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U21A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 21 0
1 U
7125 0 0
2
43495 0
0
14 Logic Display~
6 1120 196 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3641 0 0
2
43495 0
0
14 Logic Display~
6 1086 197 0 1 2
10 25
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9821 0 0
2
43495 0
0
14 Logic Display~
6 1051 199 0 1 2
10 36
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3187 0 0
2
43495 0
0
5 4071~
219 850 766 0 3 22
0 42 37 36
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U19B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 19 0
1 U
762 0 0
2
43495 0
0
8 4-In OR~
219 719 882 0 5 22
0 41 40 39 38 37
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U20B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 20 0
1 U
39 0 0
2
43495 0
0
8 4-In OR~
219 717 685 0 5 22
0 46 45 44 43 42
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U20A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 20 0
1 U
9450 0 0
2
43495 0
0
5 4071~
219 831 242 0 3 22
0 49 48 47
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 19 0
1 U
3236 0 0
2
43495 0
0
14 Logic Display~
6 1015 201 0 1 2
10 47
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3321 0 0
2
43495 0
0
8 4-In OR~
219 729 399 0 5 22
0 53 52 51 50 48
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 18 0
1 U
8879 0 0
2
43495 0
0
8 4-In OR~
219 719 155 0 5 22
0 57 56 55 54 49
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U18A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 18 0
1 U
5433 0 0
2
43495 0
0
5 4049~
219 390 2091 0 2 22
0 58 60
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U17C
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 17 0
1 U
3679 0 0
2
43495 0
0
5 4049~
219 265 2086 0 2 22
0 59 12
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U17B
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 17 0
1 U
9342 0 0
2
43495 0
0
5 4049~
219 131 2080 0 2 22
0 61 10
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U17A
17 -2 45 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 17 0
1 U
3623 0 0
2
43495 0
0
5 4082~
219 573 2014 0 5 22
0 7 61 59 58 16
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 16 0
1 U
3722 0 0
2
43495 0
0
5 4082~
219 574 1964 0 5 22
0 2 61 59 60 17
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
8993 0 0
2
43495 0
0
5 4082~
219 574 1911 0 5 22
0 3 61 12 58 18
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 15 0
1 U
3723 0 0
2
43495 0
0
5 4082~
219 573 1852 0 5 22
0 5 61 12 60 19
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 15 0
1 U
6244 0 0
2
43495 0
0
5 4082~
219 568 1789 0 5 22
0 3 10 59 58 21
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
6421 0 0
2
43495 0
0
5 4082~
219 564 1729 0 5 22
0 2 10 59 60 22
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U14A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
7743 0 0
2
43495 0
0
5 4082~
219 564 1671 0 5 22
0 8 10 10 58 23
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U13B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
9840 0 0
2
43495 0
0
5 4082~
219 561 1621 0 5 22
0 6 10 12 60 24
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U13A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
6910 0 0
2
43495 0
0
5 4082~
219 561 1496 0 5 22
0 7 61 59 58 27
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U12B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 12 0
1 U
449 0 0
2
43495 0
0
5 4082~
219 562 1444 0 5 22
0 2 61 59 60 28
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U12A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
8761 0 0
2
43495 0
0
5 4082~
219 560 1394 0 5 22
0 4 61 12 58 29
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U11B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 11 0
1 U
6748 0 0
2
43495 0
0
5 4082~
219 559 1341 0 5 22
0 6 61 12 60 30
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U11A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 11 0
1 U
7393 0 0
2
43495 0
0
5 4082~
219 557 1289 0 5 22
0 4 10 59 58 32
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
7699 0 0
2
43495 0
0
5 4082~
219 554 1232 0 5 22
0 6 10 59 62 33
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 10 0
1 U
6638 0 0
2
43495 0
0
5 4082~
219 553 1169 0 5 22
0 9 10 12 58 34
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
4595 0 0
2
43495 0
0
5 4082~
219 554 1113 0 5 22
0 3 10 12 60 35
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
9395 0 0
2
43495 0
0
5 4082~
219 551 990 0 5 22
0 7 61 59 58 38
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
3303 0 0
2
43495 0
0
5 4082~
219 548 942 0 5 22
0 2 61 59 60 39
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
4498 0 0
2
43495 0
0
5 4082~
219 550 890 0 5 22
0 5 61 12 58 40
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
9728 0 0
2
43495 0
0
5 4082~
219 547 832 0 5 22
0 3 61 12 60 41
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
3789 0 0
2
43495 0
0
5 4082~
219 544 781 0 5 22
0 5 10 59 58 43
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
3978 0 0
2
43495 0
0
5 4082~
219 543 726 0 5 22
0 3 10 59 60 44
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3494 0 0
2
43495 0
0
5 4082~
219 543 673 0 5 22
0 11 10 12 58 45
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
3507 0 0
2
43495 0
0
5 4082~
219 543 611 0 5 22
0 4 10 12 60 46
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
5151 0 0
2
43495 0
0
5 4082~
219 544 476 0 5 22
0 7 61 59 58 50
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
3701 0 0
2
43495 0
0
5 4082~
219 542 426 0 5 22
0 2 61 59 60 51
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
8585 0 0
2
43495 0
0
5 4082~
219 541 373 0 5 22
0 6 61 12 58 52
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
8809 0 0
2
43495 0
0
5 4082~
219 539 316 0 5 22
0 4 61 12 60 53
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
5993 0 0
2
43495 0
0
5 4082~
219 536 257 0 5 22
0 2 10 59 58 54
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
8654 0 0
2
43495 0
0
5 4082~
219 534 207 0 5 22
0 4 10 59 60 55
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
7223 0 0
2
43495 0
0
5 4082~
219 534 146 0 5 22
0 13 10 12 58 56
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
3641 0 0
2
43495 0
0
5 4082~
219 532 81 0 5 22
0 5 10 12 60 57
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
3104 0 0
2
43495 0
0
179
1 0 3 0 0 4096 0 35 0 0 9 3
550 1898
175 1898
175 1779
1 0 4 0 0 4096 0 43 0 0 10 3
536 1381
332 1381
332 1275
1 0 5 0 0 4096 0 51 0 0 5 2
526 877
439 877
1 0 6 0 0 4096 0 59 0 0 27 2
517 360
53 360
0 1 5 0 0 4224 0 0 36 11 0 3
439 765
439 1839
549 1839
1 0 6 0 0 4096 0 44 0 0 27 2
535 1328
53 1328
1 0 3 0 0 0 0 52 0 0 30 2
523 819
175 819
1 0 4 0 0 0 0 60 0 0 36 2
515 303
332 303
0 1 3 0 0 4096 0 0 37 30 0 4
175 1100
175 1779
544 1779
544 1776
0 1 4 0 0 4224 0 0 45 36 0 3
332 598
332 1276
533 1276
0 1 5 0 0 0 0 0 53 39 0 3
439 40
439 768
520 768
0 1 2 0 0 4096 0 0 61 24 0 3
465 413
465 244
512 244
1 0 2 0 0 0 0 38 0 0 18 2
540 1716
486 1716
1 0 6 0 0 0 0 46 0 0 27 2
530 1219
53 1219
1 0 3 0 0 0 0 54 0 0 30 2
519 713
175 713
1 0 4 0 0 0 0 62 0 0 36 2
510 194
332 194
0 0 2 0 0 4096 0 0 0 18 23 2
486 1431
486 929
1 1 2 0 0 8320 0 34 42 0 0 4
550 1951
486 1951
486 1431
538 1431
0 1 7 0 0 4224 0 0 33 20 0 3
504 1482
504 2001
549 2001
0 1 7 0 0 0 0 0 41 21 0 3
504 977
504 1483
537 1483
0 1 7 0 0 0 0 0 49 22 0 3
504 551
504 977
527 977
1 1 7 0 0 0 0 8 57 0 0 7
887 593
887 609
794 609
794 551
502 551
502 463
520 463
0 1 2 0 0 0 0 0 50 24 0 3
465 514
465 929
524 929
1 1 2 0 0 0 0 9 58 0 0 5
884 488
884 514
465 514
465 413
518 413
2 1 8 0 0 4224 0 10 39 0 0 3
101 26
101 1658
540 1658
1 1 6 0 0 0 0 7 10 0 0 3
53 50
65 50
65 26
1 1 6 0 0 4224 0 7 40 0 0 3
53 50
53 1608
537 1608
2 1 9 0 0 4224 0 11 47 0 0 3
221 25
221 1156
529 1156
0 1 3 0 0 0 0 0 11 30 0 3
175 46
185 46
185 25
1 1 3 0 0 8320 0 6 48 0 0 4
168 46
175 46
175 1100
530 1100
2 0 10 0 0 4096 0 47 0 0 176 2
529 1165
134 1165
2 1 11 0 0 4224 0 12 55 0 0 3
340 16
340 660
519 660
3 0 12 0 0 4096 0 55 0 0 170 2
519 678
268 678
2 0 10 0 0 0 0 55 0 0 176 2
519 669
134 669
0 1 4 0 0 0 0 0 12 36 0 3
301 45
304 45
304 16
1 1 4 0 0 0 0 5 56 0 0 4
294 45
332 45
332 598
519 598
2 1 13 0 0 8320 0 13 63 0 0 4
462 12
469 12
469 133
510 133
0 1 5 0 0 0 0 0 13 39 0 3
421 40
421 12
426 12
1 1 5 0 0 0 0 4 64 0 0 4
401 40
477 40
477 68
508 68
1 3 14 0 0 4224 0 20 16 0 0 3
1120 214
1120 1796
959 1796
5 2 15 0 0 8320 0 14 16 0 0 4
770 1921
855 1921
855 1805
913 1805
5 4 16 0 0 4224 0 33 14 0 0 4
594 2014
686 2014
686 1935
720 1935
5 3 17 0 0 4224 0 34 14 0 0 4
595 1964
662 1964
662 1926
720 1926
5 2 18 0 0 12416 0 35 14 0 0 4
595 1911
630 1911
630 1917
720 1917
5 1 19 0 0 12416 0 36 14 0 0 4
594 1852
646 1852
646 1908
720 1908
5 1 20 0 0 8320 0 15 16 0 0 4
762 1670
846 1670
846 1787
913 1787
5 4 21 0 0 8320 0 37 15 0 0 4
589 1789
644 1789
644 1684
712 1684
5 3 22 0 0 12416 0 38 15 0 0 4
585 1729
615 1729
615 1675
712 1675
5 2 23 0 0 4224 0 39 15 0 0 4
585 1671
692 1671
692 1666
712 1666
1 5 24 0 0 12416 0 15 40 0 0 4
712 1657
649 1657
649 1621
582 1621
1 3 25 0 0 4224 0 21 17 0 0 3
1086 215
1086 1276
925 1276
5 2 26 0 0 4224 0 18 17 0 0 3
778 1405
778 1285
879 1285
5 4 27 0 0 12416 0 41 18 0 0 4
582 1496
636 1496
636 1419
728 1419
5 3 28 0 0 12416 0 42 18 0 0 4
583 1444
611 1444
611 1410
728 1410
5 2 29 0 0 12416 0 43 18 0 0 4
581 1394
630 1394
630 1401
728 1401
5 1 30 0 0 4224 0 44 18 0 0 4
580 1341
675 1341
675 1392
728 1392
5 1 31 0 0 8320 0 19 17 0 0 4
775 1181
832 1181
832 1267
879 1267
5 4 32 0 0 8320 0 45 19 0 0 4
578 1289
671 1289
671 1195
725 1195
5 3 33 0 0 12416 0 46 19 0 0 4
575 1232
640 1232
640 1186
725 1186
5 2 34 0 0 4224 0 47 19 0 0 4
574 1169
680 1169
680 1177
725 1177
5 1 35 0 0 4224 0 48 19 0 0 4
575 1113
709 1113
709 1168
725 1168
3 1 36 0 0 8320 0 23 22 0 0 3
883 766
1051 766
1051 217
5 2 37 0 0 4224 0 24 23 0 0 3
752 882
752 775
837 775
5 4 38 0 0 8320 0 49 24 0 0 4
572 990
657 990
657 896
702 896
5 3 39 0 0 20608 0 50 24 0 0 6
569 942
622 942
622 899
627 899
627 887
702 887
5 2 40 0 0 12416 0 51 24 0 0 4
571 890
620 890
620 878
702 878
5 1 41 0 0 4224 0 52 24 0 0 4
568 832
689 832
689 869
702 869
5 1 42 0 0 8320 0 25 23 0 0 4
750 685
779 685
779 757
837 757
5 4 43 0 0 4224 0 53 25 0 0 4
565 781
654 781
654 699
700 699
5 3 44 0 0 12416 0 54 25 0 0 4
564 726
627 726
627 690
700 690
5 2 45 0 0 4224 0 55 25 0 0 4
564 673
637 673
637 681
700 681
5 1 46 0 0 4224 0 56 25 0 0 4
564 611
680 611
680 672
700 672
3 1 47 0 0 4224 0 26 27 0 0 3
864 242
1015 242
1015 219
5 2 48 0 0 8320 0 28 26 0 0 4
762 399
791 399
791 251
818 251
5 1 49 0 0 4224 0 29 26 0 0 3
752 155
752 233
818 233
5 4 50 0 0 4224 0 57 28 0 0 4
565 476
647 476
647 413
712 413
5 3 51 0 0 12416 0 58 28 0 0 4
563 426
624 426
624 404
712 404
5 2 52 0 0 12416 0 59 28 0 0 4
562 373
634 373
634 395
712 395
5 1 53 0 0 4224 0 60 28 0 0 4
560 316
670 316
670 386
712 386
5 4 54 0 0 4224 0 61 29 0 0 4
557 257
687 257
687 169
702 169
5 3 55 0 0 4224 0 62 29 0 0 4
555 207
656 207
656 160
702 160
5 2 56 0 0 4224 0 63 29 0 0 4
555 146
681 146
681 151
702 151
5 1 57 0 0 4224 0 64 29 0 0 4
553 81
696 81
696 142
702 142
4 0 58 0 0 4096 0 33 0 0 162 2
549 2028
366 2028
3 0 59 0 0 4096 0 33 0 0 154 2
549 2019
234 2019
4 0 60 0 0 4096 0 34 0 0 168 2
550 1978
393 1978
3 0 59 0 0 4096 0 34 0 0 154 2
550 1969
234 1969
4 0 58 0 0 4096 0 35 0 0 162 2
550 1925
366 1925
3 0 12 0 0 4096 0 35 0 0 172 2
550 1916
268 1916
4 0 60 0 0 0 0 36 0 0 168 2
549 1866
393 1866
3 0 12 0 0 0 0 36 0 0 172 2
549 1857
268 1857
4 0 58 0 0 0 0 41 0 0 161 2
537 1510
366 1510
3 0 59 0 0 0 0 41 0 0 152 2
537 1501
234 1501
4 0 60 0 0 0 0 42 0 0 167 2
538 1458
393 1458
3 0 59 0 0 0 0 42 0 0 152 2
538 1449
234 1449
4 0 58 0 0 0 0 43 0 0 161 2
536 1408
366 1408
3 0 12 0 0 0 0 43 0 0 171 2
536 1399
268 1399
4 0 60 0 0 0 0 44 0 0 167 2
535 1355
393 1355
3 0 12 0 0 0 0 44 0 0 171 2
535 1346
268 1346
4 0 58 0 0 0 0 49 0 0 159 2
527 1004
366 1004
3 0 59 0 0 0 0 49 0 0 151 2
527 995
234 995
4 0 60 0 0 0 0 50 0 0 166 2
524 956
393 956
3 0 59 0 0 0 0 50 0 0 151 2
524 947
234 947
4 0 58 0 0 0 0 51 0 0 159 2
526 904
366 904
3 0 12 0 0 0 0 51 0 0 170 2
526 895
268 895
4 0 60 0 0 0 0 52 0 0 166 2
523 846
393 846
3 0 12 0 0 0 0 52 0 0 170 2
523 837
268 837
4 0 58 0 0 0 0 57 0 0 158 2
520 490
366 490
3 0 59 0 0 0 0 57 0 0 150 2
520 481
234 481
4 0 60 0 0 0 0 58 0 0 165 2
518 440
393 440
3 0 59 0 0 0 0 58 0 0 150 2
518 431
234 431
4 0 58 0 0 0 0 59 0 0 158 2
517 387
366 387
3 0 12 0 0 0 0 59 0 0 169 2
517 378
268 378
4 0 60 0 0 0 0 60 0 0 165 2
515 330
393 330
3 0 12 0 0 0 0 60 0 0 169 2
515 321
268 321
2 0 61 0 0 4096 0 57 0 0 119 2
520 472
106 472
2 0 61 0 0 0 0 58 0 0 119 2
518 422
106 422
2 0 61 0 0 0 0 59 0 0 119 2
517 369
106 369
0 2 61 0 0 4224 0 0 60 122 0 3
106 828
106 312
515 312
2 0 61 0 0 0 0 50 0 0 122 2
524 938
106 938
2 0 61 0 0 0 0 51 0 0 122 2
526 886
106 886
0 2 61 0 0 0 0 0 52 123 0 3
106 989
106 828
523 828
0 2 61 0 0 0 0 0 49 127 0 3
106 1340
106 986
527 986
2 0 61 0 0 0 0 41 0 0 127 2
537 1492
106 1492
2 0 61 0 0 0 0 42 0 0 127 2
538 1440
106 1440
2 0 61 0 0 0 0 43 0 0 127 2
536 1390
106 1390
0 2 61 0 0 0 0 0 44 131 0 3
106 1848
106 1337
535 1337
2 0 61 0 0 0 0 33 0 0 131 2
549 2010
106 2010
2 0 61 0 0 0 0 34 0 0 131 2
550 1960
106 1960
2 0 61 0 0 0 0 35 0 0 131 2
550 1907
106 1907
0 2 61 0 0 0 0 0 36 179 0 3
106 2116
106 1848
549 1848
4 0 58 0 0 0 0 37 0 0 162 2
544 1803
366 1803
3 0 59 0 0 0 0 37 0 0 154 2
544 1794
234 1794
2 0 10 0 0 4096 0 37 0 0 176 2
544 1785
134 1785
4 0 58 0 0 0 0 45 0 0 161 2
533 1303
366 1303
3 0 59 0 0 0 0 45 0 0 152 2
533 1294
234 1294
2 0 10 0 0 0 0 45 0 0 176 2
533 1285
134 1285
0 0 60 0 0 0 0 0 0 0 167 2
534 1249
393 1249
2 0 10 0 0 0 0 46 0 0 176 2
530 1228
134 1228
4 0 58 0 0 0 0 53 0 0 159 2
520 795
366 795
3 0 59 0 0 0 0 53 0 0 151 2
520 786
234 786
2 0 10 0 0 0 0 53 0 0 176 2
520 777
134 777
4 0 58 0 0 0 0 61 0 0 158 2
512 271
366 271
3 0 59 0 0 0 0 61 0 0 150 2
512 262
234 262
2 0 10 0 0 0 0 61 0 0 176 2
512 253
134 253
4 0 60 0 0 0 0 54 0 0 166 2
519 740
393 740
2 0 10 0 0 0 0 54 0 0 176 2
519 722
134 722
4 0 60 0 0 0 0 62 0 0 165 2
510 221
393 221
2 0 10 0 0 0 0 62 0 0 176 2
510 203
134 203
0 3 59 0 0 4224 0 0 62 151 0 3
234 734
234 212
510 212
0 3 59 0 0 0 0 0 54 152 0 3
234 1239
234 731
519 731
0 3 59 0 0 0 0 0 46 154 0 3
234 1735
234 1237
530 1237
0 4 60 0 0 0 0 0 38 168 0 3
393 1742
393 1743
540 1743
0 3 59 0 0 0 0 0 38 178 0 3
234 2111
234 1734
540 1734
2 0 10 0 0 0 0 38 0 0 176 2
540 1725
134 1725
3 0 12 0 0 0 0 63 0 0 169 2
510 151
268 151
2 0 10 0 0 0 0 63 0 0 176 2
510 142
134 142
0 4 58 0 0 4224 0 0 63 159 0 3
366 687
366 160
510 160
0 4 58 0 0 0 0 0 55 161 0 3
366 1184
366 687
519 687
0 3 12 0 0 0 0 0 47 171 0 2
268 1174
529 1174
0 4 58 0 0 0 0 0 47 162 0 3
366 1687
366 1183
529 1183
0 4 58 0 0 0 0 0 39 177 0 3
366 2102
366 1685
540 1685
3 0 10 0 0 0 0 39 0 0 176 2
540 1676
134 1676
2 0 10 0 0 0 0 39 0 0 176 2
540 1667
134 1667
0 4 60 0 0 4224 0 0 64 166 0 3
393 625
393 95
508 95
0 4 60 0 0 0 0 0 56 167 0 3
393 1130
393 625
519 625
0 4 60 0 0 0 0 0 48 168 0 3
393 1639
393 1127
530 1127
2 4 60 0 0 0 0 30 40 0 0 3
393 2073
393 1635
537 1635
0 3 12 0 0 4224 0 0 64 170 0 3
268 617
268 86
508 86
0 3 12 0 0 0 0 0 56 171 0 3
268 1120
268 616
519 616
0 3 12 0 0 0 0 0 48 172 0 3
268 1629
268 1118
530 1118
2 3 12 0 0 0 0 31 40 0 0 3
268 2068
268 1626
537 1626
0 2 10 0 0 0 0 0 40 176 0 3
134 1615
134 1617
537 1617
0 2 10 0 0 0 0 0 48 176 0 3
134 1106
134 1109
530 1109
0 2 10 0 0 0 0 0 56 176 0 3
134 609
134 607
519 607
2 2 10 0 0 4224 0 32 64 0 0 3
134 2062
134 77
508 77
1 1 58 0 0 0 0 1 30 0 0 5
346 2102
367 2102
367 2112
393 2112
393 2109
1 1 59 0 0 0 0 2 31 0 0 3
214 2111
268 2111
268 2104
1 1 61 0 0 0 0 3 32 0 0 3
87 2116
134 2116
134 2098
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
