CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
42
13 Logic Switch~
5 102 376 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 b2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4139 0 0
2
5.89884e-315 0
0
13 Logic Switch~
5 111 272 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 a2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6435 0 0
2
5.89884e-315 5.26354e-315
0
13 Logic Switch~
5 228 383 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 b1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5283 0 0
2
5.89884e-315 5.30499e-315
0
13 Logic Switch~
5 229 284 0 1 11
0 39
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 a1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6874 0 0
2
5.89884e-315 5.32571e-315
0
13 Logic Switch~
5 298 77 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5305 0 0
2
5.89884e-315 5.34643e-315
0
13 Logic Switch~
5 224 79 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 s0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
5.89884e-315 5.3568e-315
0
13 Logic Switch~
5 134 78 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 s1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
969 0 0
2
5.89884e-315 5.36716e-315
0
5 4049~
219 152 1053 0 2 22
0 3 2
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 2 0
1 U
8402 0 0
2
43537.2 0
0
14 Logic Display~
6 931 100 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
43537.2 0
0
5 4071~
219 1084 1204 0 3 22
0 5 6 4
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
4292 0 0
2
43537.2 0
0
5 4081~
219 1007 1280 0 3 22
0 8 7 6
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
6118 0 0
2
43537.2 0
0
5 4030~
219 930 1258 0 3 22
0 10 9 8
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U9B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
34 0 0
2
43537.2 0
0
5 4081~
219 929 1184 0 3 22
0 10 9 5
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
6357 0 0
2
43537.2 0
0
14 Logic Display~
6 1070 107 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
319 0 0
2
43537.2 0
0
5 4030~
219 1016 998 0 3 22
0 12 7 11
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U9A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
3976 0 0
2
43537.2 0
0
5 4030~
219 929 958 0 3 22
0 10 9 12
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
7634 0 0
2
43537.2 0
0
5 4071~
219 803 1094 0 3 22
0 14 13 9
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
523 0 0
2
43537.2 0
0
5 4081~
219 731 1146 0 3 22
0 15 3 13
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
6748 0 0
2
43537.2 0
0
5 4073~
219 731 1067 0 4 22
0 17 16 2 14
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U8A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 8 0
1 U
6901 0 0
2
43537.2 0
0
5 4071~
219 817 919 0 3 22
0 19 18 10
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
842 0 0
2
43537.2 0
0
5 4049~
219 386 911 0 2 22
0 21 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 2 0
1 U
3277 0 0
2
43537.2 0
0
5 4073~
219 737 972 0 4 22
0 15 22 20 18
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 4 0
1 U
4212 0 0
2
43537.2 0
0
5 4081~
219 737 887 0 3 22
0 23 21 19
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
4720 0 0
2
43537.2 0
0
5 4071~
219 654 861 0 3 22
0 17 16 23
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 18
65 0 0 0 4 1 7 0
1 U
5551 0 0
2
43537.2 0
0
5 4071~
219 1020 661 0 3 22
0 26 25 7
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
6986 0 0
2
43537.2 1
0
5 4081~
219 877 692 0 3 22
0 28 27 25
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
8745 0 0
2
43537.2 2
0
5 4081~
219 961 613 0 3 22
0 29 24 26
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
9592 0 0
2
43537.2 3
0
5 4030~
219 870 604 0 3 22
0 28 27 29
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8748 0 0
2
43537.2 4
0
14 Logic Display~
6 1134 107 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7168 0 0
2
43537.2 5
0
5 4030~
219 897 372 0 3 22
0 31 24 30
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
631 0 0
2
43537.2 6
0
5 4030~
219 819 307 0 3 22
0 28 27 31
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
9466 0 0
2
43537.2 7
0
5 4071~
219 706 411 0 3 22
0 33 32 27
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3266 0 0
2
43537.2 8
0
5 4081~
219 623 451 0 3 22
0 15 34 32
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
7693 0 0
2
43537.2 9
0
5 4049~
219 297 399 0 2 22
0 34 35
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 2 0
1 U
3723 0 0
2
43537.2 10
0
5 4073~
219 622 387 0 4 22
0 17 15 35 33
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 4 0
1 U
3440 0 0
2
43537.2 11
0
5 4071~
219 719 251 0 3 22
0 37 36 28
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
6263 0 0
2
43537.2 12
0
5 4049~
219 284 328 0 2 22
0 39 38
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 2 0
1 U
4900 0 0
2
43537.2 13
0
5 4049~
219 276 137 0 2 22
0 16 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 2 0
1 U
8783 0 0
2
43537.2 14
0
5 4073~
219 622 311 0 4 22
0 15 22 38 36
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
3221 0 0
2
43537.2 15
0
5 4081~
219 620 224 0 3 22
0 40 39 37
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3215 0 0
2
43537.2 16
0
5 4049~
219 174 137 0 2 22
0 15 17
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U2A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 2 0
1 U
7903 0 0
2
43537.2 17
0
5 4071~
219 520 207 0 3 22
0 16 17 40
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
7121 0 0
2
43537.2 18
0
65
2 3 2 0 0 12416 0 8 19 0 0 4
173 1053
193 1053
193 1076
707 1076
1 0 3 0 0 0 0 8 0 0 20 2
137 1053
137 1053
1 3 4 0 0 16512 0 9 10 0 0 6
931 118
983 118
983 151
1198 151
1198 1204
1117 1204
3 1 5 0 0 12416 0 13 10 0 0 4
950 1184
973 1184
973 1195
1071 1195
3 2 6 0 0 8320 0 11 10 0 0 4
1028 1280
1053 1280
1053 1213
1071 1213
0 2 7 0 0 20480 0 0 11 13 0 6
991 1003
903 1003
903 1124
813 1124
813 1289
983 1289
3 1 8 0 0 8320 0 12 11 0 0 4
963 1258
971 1258
971 1271
983 1271
0 2 9 0 0 4096 0 0 12 10 0 3
861 1193
861 1267
914 1267
0 1 10 0 0 4096 0 0 12 11 0 3
873 1175
873 1249
914 1249
0 2 9 0 0 4096 0 0 13 15 0 3
846 1094
846 1193
905 1193
0 1 10 0 0 4224 0 0 13 16 0 3
859 948
859 1175
905 1175
1 3 11 0 0 12416 0 14 15 0 0 5
1070 125
1070 466
1149 466
1149 998
1049 998
3 2 7 0 0 8320 0 25 15 0 0 6
1053 661
1063 661
1063 946
991 946
991 1007
1000 1007
3 1 12 0 0 16512 0 16 15 0 0 5
962 958
962 977
978 977
978 989
1000 989
3 2 9 0 0 8320 0 17 16 0 0 4
836 1094
872 1094
872 967
913 967
3 1 10 0 0 0 0 20 16 0 0 4
850 919
859 919
859 949
913 949
3 2 13 0 0 8320 0 18 17 0 0 4
752 1146
782 1146
782 1103
790 1103
4 1 14 0 0 12416 0 19 17 0 0 4
752 1067
766 1067
766 1085
790 1085
0 1 15 0 0 8192 0 0 18 28 0 3
166 963
166 1137
707 1137
1 2 3 0 0 28800 0 1 18 0 0 8
114 376
130 376
130 411
79 411
79 909
137 909
137 1155
707 1155
0 2 16 0 0 8192 0 0 19 31 0 3
348 870
348 1067
707 1067
1 0 17 0 0 4096 0 19 0 0 32 3
707 1058
268 1058
268 852
4 2 18 0 0 8320 0 22 20 0 0 4
758 972
773 972
773 928
804 928
3 1 19 0 0 12416 0 23 20 0 0 4
758 887
778 887
778 910
804 910
2 3 20 0 0 4224 0 21 22 0 0 4
407 911
572 911
572 981
713 981
0 1 21 0 0 4096 0 0 21 29 0 3
366 896
366 911
371 911
0 2 22 0 0 4224 0 0 22 58 0 3
321 311
321 972
713 972
0 1 15 0 0 12416 0 0 22 64 0 5
146 136
146 239
166 239
166 963
713 963
1 2 21 0 0 8320 0 2 23 0 0 4
123 272
147 272
147 896
713 896
3 1 23 0 0 4224 0 24 23 0 0 4
687 861
704 861
704 878
713 878
0 2 16 0 0 4224 0 0 24 65 0 3
327 198
327 870
641 870
0 1 17 0 0 4224 0 0 24 63 0 3
199 137
199 852
641 852
0 2 24 0 0 8192 0 0 27 34 0 3
547 489
547 622
937 622
1 2 24 0 0 8320 0 5 30 0 0 6
310 77
432 77
432 489
819 489
819 381
881 381
3 2 25 0 0 4224 0 26 25 0 0 4
898 692
967 692
967 670
1007 670
3 1 26 0 0 4224 0 27 25 0 0 3
982 613
982 652
1007 652
0 2 27 0 0 4096 0 0 26 40 0 3
769 613
769 701
853 701
0 1 28 0 0 8192 0 0 26 41 0 3
758 594
758 683
853 683
1 3 29 0 0 4224 0 27 28 0 0 2
937 604
903 604
0 2 27 0 0 4224 0 0 28 44 0 3
769 411
769 613
854 613
0 1 28 0 0 4224 0 0 28 45 0 3
758 251
758 595
854 595
3 1 30 0 0 8320 0 30 29 0 0 3
930 372
1134 372
1134 125
3 1 31 0 0 8320 0 31 30 0 0 4
852 307
866 307
866 363
881 363
3 2 27 0 0 0 0 32 31 0 0 4
739 411
772 411
772 316
803 316
3 1 28 0 0 0 0 36 31 0 0 4
752 251
774 251
774 298
803 298
3 2 32 0 0 8320 0 33 32 0 0 4
644 451
667 451
667 420
693 420
4 1 33 0 0 12416 0 35 32 0 0 4
643 387
667 387
667 402
693 402
0 2 34 0 0 8320 0 0 33 51 0 3
260 383
260 460
599 460
0 1 15 0 0 128 0 0 33 52 0 3
341 387
341 442
599 442
2 3 35 0 0 4224 0 34 35 0 0 4
318 399
578 399
578 396
598 396
1 1 34 0 0 0 0 3 34 0 0 4
240 383
274 383
274 399
282 399
0 2 15 0 0 0 0 0 35 60 0 3
341 302
341 387
598 387
0 1 17 0 0 0 0 0 35 63 0 3
395 216
395 378
598 378
4 2 36 0 0 8320 0 39 36 0 0 4
643 311
680 311
680 260
706 260
3 1 37 0 0 12416 0 40 36 0 0 4
641 224
671 224
671 242
706 242
2 3 38 0 0 12416 0 37 39 0 0 4
305 328
437 328
437 320
598 320
0 1 39 0 0 4096 0 0 37 61 0 3
261 284
261 328
269 328
2 2 22 0 0 128 0 38 39 0 0 3
297 137
297 311
598 311
1 0 16 0 0 0 0 38 0 0 65 2
261 137
236 137
0 1 15 0 0 0 0 0 39 64 0 4
146 111
341 111
341 302
598 302
1 2 39 0 0 4224 0 4 40 0 0 4
241 284
503 284
503 233
596 233
3 1 40 0 0 12416 0 42 40 0 0 4
553 207
567 207
567 215
596 215
2 2 17 0 0 128 0 41 42 0 0 4
195 137
225 137
225 216
507 216
1 1 15 0 0 0 0 7 41 0 0 3
146 78
146 137
159 137
1 1 16 0 0 128 0 6 42 0 0 3
236 79
236 198
507 198
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
