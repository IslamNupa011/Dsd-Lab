CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
66
13 Logic Switch~
5 193 32 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43493.3 0
0
13 Logic Switch~
5 285 29 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
43493.3 1
0
13 Logic Switch~
5 490 2451 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
43493.3 2
0
13 Logic Switch~
5 637 2441 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 s1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43493.3 3
0
13 Logic Switch~
5 778 2436 0 1 11
0 33
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
43493.3 4
0
13 Logic Switch~
5 30 40 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.89879e-315 0
0
13 Logic Switch~
5 122 37 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89879e-315 5.26354e-315
0
5 4049~
219 242 127 0 2 22
0 3 8
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U15C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 15 0
1 U
7361 0 0
2
43493.3 5
0
5 4049~
219 320 126 0 2 22
0 6 7
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U15D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 15 0
1 U
4747 0 0
2
43493.3 6
0
14 Logic Display~
6 1461 240 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
43493.3 7
0
14 Logic Display~
6 1424 244 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
43493.3 8
0
2 +V
167 1289 2351 0 1 3
0 11
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
43493.3 9
0
7 Ground~
168 1268 1820 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
43493.3 10
0
5 4082~
219 1040 1313 0 5 22
0 3 38 37 36 32
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U23B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 23 0
1 U
4597 0 0
2
43493.3 11
0
5 4082~
219 1042 1380 0 5 22
0 8 38 37 33 31
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U23A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 23 0
1 U
3835 0 0
2
43493.3 12
0
5 4082~
219 1044 1444 0 5 22
0 4 38 34 36 30
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U22B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 22 0
1 U
3670 0 0
2
43493.3 13
0
5 4082~
219 1046 1507 0 5 22
0 6 38 34 33 29
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U22A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 22 0
1 U
5616 0 0
2
43493.3 14
0
5 4082~
219 1048 1565 0 5 22
0 4 35 37 36 65
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U21B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 2 21 0
1 U
9323 0 0
2
43493.3 15
0
5 4082~
219 1048 1631 0 5 22
0 6 35 37 33 27
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U21A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 21 0
1 U
317 0 0
2
43493.3 16
0
5 4082~
219 1049 1691 0 5 22
0 2 35 34 36 26
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U20B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 20 0
1 U
3108 0 0
2
43493.3 17
0
5 4082~
219 1050 1746 0 5 22
0 11 35 34 33 25
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U20A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 20 0
1 U
4299 0 0
2
43493.3 18
0
5 4082~
219 1048 1908 0 5 22
0 6 38 37 36 22
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U19B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 19 0
1 U
9672 0 0
2
43493.3 19
0
5 4082~
219 1048 1968 0 5 22
0 7 38 37 33 21
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U19A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 19 0
1 U
7876 0 0
2
43493.3 20
0
5 4082~
219 1048 2025 0 5 22
0 3 38 34 36 20
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U18B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 18 0
1 U
6369 0 0
2
43493.3 21
0
5 4082~
219 1048 2087 0 5 22
0 2 38 34 33 19
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U18A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 18 0
1 U
9172 0 0
2
43493.3 22
0
5 4082~
219 1050 2144 0 5 22
0 3 35 37 36 18
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U17B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 17 0
1 U
7100 0 0
2
43493.3 23
0
5 4082~
219 1052 2200 0 5 22
0 5 35 37 33 17
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U17A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 17 0
1 U
3820 0 0
2
43493.3 24
0
5 4082~
219 1052 2256 0 5 22
0 2 35 34 36 16
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 16 0
1 U
7678 0 0
2
43493.3 25
0
5 4082~
219 1053 2312 0 5 22
0 11 35 34 33 15
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U16A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
961 0 0
2
43493.3 26
0
5 4049~
219 541 2421 0 2 22
0 35 38
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U15B
13 -2 41 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 15 0
1 U
3178 0 0
2
43493.3 27
0
5 4049~
219 696 2418 0 2 22
0 34 37
0
0 0 624 90
4 4049
-7 -24 21 -16
4 U15A
13 -2 41 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 15 0
1 U
3409 0 0
2
43493.3 28
0
5 4049~
219 841 2413 0 2 22
0 33 36
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U1F
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 1 0
1 U
3951 0 0
2
43493.3 29
0
8 4-In OR~
219 1152 1414 0 5 22
0 32 31 30 29 24
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U14B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 14 0
1 U
8885 0 0
2
43493.3 30
0
8 4-In OR~
219 1157 1614 0 5 22
0 28 27 26 25 23
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U14A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 14 0
1 U
3780 0 0
2
43493.3 31
0
5 4071~
219 1234 1484 0 3 22
0 24 23 10
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
9265 0 0
2
43493.3 32
0
8 4-In OR~
219 1168 2018 0 5 22
0 22 21 20 19 12
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U13B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
9442 0 0
2
43493.3 33
0
8 4-In OR~
219 1176 2214 0 5 22
0 18 17 16 15 13
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U13A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
9424 0 0
2
43493.3 34
0
5 4071~
219 1292 2034 0 3 22
0 12 13 9
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
9968 0 0
2
43493.3 35
0
14 Logic Display~
6 1385 247 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
43493.3 36
0
5 4071~
219 1280 822 0 3 22
0 43 44 39
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
8464 0 0
2
5.89879e-315 5.30499e-315
0
8 4-In OR~
219 1164 1002 0 5 22
0 49 48 47 46 44
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 12 0
1 U
7168 0 0
2
5.89879e-315 5.32571e-315
0
8 4-In OR~
219 1156 806 0 5 22
0 53 52 51 50 43
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
3171 0 0
2
5.89879e-315 5.34643e-315
0
14 Logic Display~
6 1345 248 0 1 2
10 54
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4139 0 0
2
5.89879e-315 5.3568e-315
0
5 4071~
219 1222 272 0 3 22
0 56 55 54
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
6435 0 0
2
5.89879e-315 5.36716e-315
0
8 4-In OR~
219 1145 402 0 5 22
0 60 59 58 57 55
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
5283 0 0
2
5.89879e-315 5.37752e-315
0
8 4-In OR~
219 1140 202 0 5 22
0 64 63 62 61 56
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
6874 0 0
2
5.89879e-315 5.38788e-315
0
5 4082~
219 1041 1100 0 5 22
0 40 35 34 33 46
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
5305 0 0
2
5.89879e-315 5.39306e-315
0
5 4082~
219 1040 1044 0 5 22
0 2 35 34 36 47
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U9A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
34 0 0
2
5.89879e-315 5.39824e-315
0
5 4082~
219 1040 988 0 5 22
0 3 35 37 33 48
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
969 0 0
2
5.89879e-315 5.40342e-315
0
5 4082~
219 1038 932 0 5 22
0 5 35 37 36 49
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
8402 0 0
2
5.89879e-315 5.4086e-315
0
5 4082~
219 1036 875 0 5 22
0 3 38 34 33 50
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
3751 0 0
2
5.89879e-315 5.41378e-315
0
5 4082~
219 1036 813 0 5 22
0 5 38 34 36 51
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
4292 0 0
2
5.89879e-315 5.41896e-315
0
5 4082~
219 1036 756 0 5 22
0 41 38 37 33 52
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
6118 0 0
2
5.89879e-315 5.42414e-315
0
5 4082~
219 1036 696 0 5 22
0 4 38 37 36 53
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
34 0 0
2
5.89879e-315 5.42933e-315
0
5 4082~
219 1038 534 0 5 22
0 40 35 34 33 57
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
6357 0 0
2
5.89879e-315 5.43192e-315
0
5 4082~
219 1037 479 0 5 22
0 2 35 34 36 58
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
319 0 0
2
5.89879e-315 5.43451e-315
0
5 4082~
219 1036 419 0 5 22
0 4 35 37 33 59
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
3976 0 0
2
5.89879e-315 5.4371e-315
0
5 4082~
219 1036 353 0 5 22
0 6 35 37 36 66
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 512 2 1 4 0
1 U
7634 0 0
2
5.89879e-315 5.43969e-315
0
5 4082~
219 1034 295 0 5 22
0 4 38 34 33 61
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
523 0 0
2
5.89879e-315 5.44228e-315
0
5 4082~
219 1032 232 0 5 22
0 2 38 34 36 62
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
6748 0 0
2
5.89879e-315 5.44487e-315
0
5 4082~
219 1030 168 0 5 22
0 42 38 37 33 63
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
6901 0 0
2
5.89879e-315 5.44746e-315
0
5 4082~
219 1028 101 0 5 22
0 5 38 37 36 64
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
842 0 0
2
5.89879e-315 5.45005e-315
0
5 4049~
219 78 117 0 2 22
0 5 42
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
3277 0 0
2
5.89879e-315 5.45264e-315
0
5 4049~
219 157 134 0 2 22
0 4 41
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U1A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
4212 0 0
2
5.89879e-315 5.45523e-315
0
7 Ground~
168 1256 608 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4720 0 0
2
5.89879e-315 5.45782e-315
0
2 +V
167 1277 1139 0 1 3
0 40
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5551 0 0
2
5.89879e-315 5.46041e-315
0
181
1 0 3 0 0 4096 0 26 0 0 13 3
1026 2131
205 2131
205 2009
1 0 4 0 0 4224 0 18 0 0 14 3
1024 1552
134 1552
134 1434
1 0 5 0 0 4096 0 50 0 0 8 2
1014 919
51 919
1 0 6 0 0 4096 0 58 0 0 21 2
1012 340
297 340
1 0 6 0 0 4096 0 19 0 0 21 2
1024 1618
297 1618
1 0 3 0 0 0 0 49 0 0 22 2
1016 975
205 975
1 0 4 0 0 0 0 57 0 0 110 2
1012 406
134 406
0 1 5 0 0 4224 0 0 27 15 0 3
51 799
51 2187
1028 2187
1 0 6 0 0 0 0 17 0 0 21 2
1022 1494
297 1494
0 1 3 0 0 0 0 0 51 22 0 4
205 866
1003 866
1003 862
1012 862
1 0 4 0 0 0 0 59 0 0 110 2
1010 282
134 282
1 0 2 0 0 4096 0 25 0 0 27 2
1024 2074
916 2074
0 1 3 0 0 0 0 0 24 22 0 3
205 1300
205 2012
1024 2012
0 1 4 0 0 128 0 0 16 110 0 4
134 681
134 1434
1020 1434
1020 1431
0 1 5 0 0 0 0 0 52 111 0 3
51 89
51 800
1012 800
0 1 2 0 0 12416 0 0 60 104 0 4
904 600
466 600
466 219
1008 219
2 1 7 0 0 4224 0 9 23 0 0 3
341 126
341 1955
1024 1955
0 1 6 0 0 0 0 0 9 21 0 3
297 124
297 126
305 126
2 1 8 0 0 4224 0 8 15 0 0 3
263 127
263 1367
1018 1367
0 1 3 0 0 0 0 0 8 22 0 3
205 126
205 127
227 127
1 1 6 0 0 4224 0 2 22 0 0 3
297 29
297 1895
1024 1895
1 1 3 0 0 4224 0 1 14 0 0 3
205 32
205 1300
1016 1300
1 3 9 0 0 4224 0 10 38 0 0 3
1461 258
1461 2034
1325 2034
1 3 10 0 0 4224 0 11 35 0 0 5
1424 262
1424 1196
1296 1196
1296 1484
1267 1484
0 1 11 0 0 4224 0 0 21 26 0 3
938 2299
938 1733
1026 1733
1 1 11 0 0 0 0 12 29 0 0 5
1289 2360
1289 2375
935 2375
935 2299
1029 2299
1 0 2 0 0 0 0 28 0 0 28 3
1028 2243
916 2243
916 1810
1 1 2 0 0 0 0 20 13 0 0 5
1025 1678
916 1678
916 1810
1268 1810
1268 1814
5 1 12 0 0 4224 0 36 38 0 0 4
1201 2018
1248 2018
1248 2025
1279 2025
5 2 13 0 0 8320 0 37 38 0 0 4
1209 2214
1251 2214
1251 2043
1279 2043
0 0 14 0 0 8320 0 0 0 0 0 3
1287 2092
1287 2093
1284 2093
5 4 15 0 0 4224 0 29 37 0 0 3
1074 2312
1159 2312
1159 2228
5 3 16 0 0 4224 0 28 37 0 0 4
1073 2256
1122 2256
1122 2219
1159 2219
5 2 17 0 0 12416 0 27 37 0 0 4
1073 2200
1089 2200
1089 2210
1159 2210
5 1 18 0 0 8320 0 26 37 0 0 4
1071 2144
1120 2144
1120 2201
1159 2201
5 4 19 0 0 8320 0 25 36 0 0 4
1069 2087
1114 2087
1114 2032
1151 2032
5 3 20 0 0 4224 0 24 36 0 0 4
1069 2025
1134 2025
1134 2023
1151 2023
5 2 21 0 0 12416 0 23 36 0 0 4
1069 1968
1094 1968
1094 2014
1151 2014
5 1 22 0 0 8320 0 22 36 0 0 4
1069 1908
1107 1908
1107 2005
1151 2005
5 2 23 0 0 8320 0 34 35 0 0 4
1190 1614
1197 1614
1197 1493
1221 1493
5 1 24 0 0 8320 0 33 35 0 0 4
1185 1414
1202 1414
1202 1475
1221 1475
5 4 25 0 0 8320 0 21 34 0 0 6
1071 1746
1101 1746
1101 1651
1113 1651
1113 1628
1140 1628
5 3 26 0 0 4224 0 20 34 0 0 5
1070 1691
1070 1638
1098 1638
1098 1619
1140 1619
5 2 27 0 0 12416 0 19 34 0 0 4
1069 1631
1088 1631
1088 1610
1140 1610
0 1 28 0 0 4224 0 0 34 0 0 4
1072 1566
1120 1566
1120 1601
1140 1601
5 4 29 0 0 8320 0 17 33 0 0 4
1067 1507
1094 1507
1094 1428
1135 1428
5 3 30 0 0 12416 0 16 33 0 0 4
1065 1444
1078 1444
1078 1419
1135 1419
5 2 31 0 0 12416 0 15 33 0 0 4
1063 1380
1094 1380
1094 1410
1135 1410
5 1 32 0 0 8320 0 14 33 0 0 4
1061 1313
1108 1313
1108 1401
1135 1401
0 4 33 0 0 4096 0 0 21 68 0 4
806 1770
1019 1770
1019 1760
1026 1760
0 3 34 0 0 4096 0 0 21 66 0 4
668 1760
1014 1760
1014 1751
1026 1751
0 2 35 0 0 4096 0 0 21 61 0 4
516 1750
1004 1750
1004 1742
1026 1742
0 4 36 0 0 8192 0 0 20 92 0 3
844 1706
844 1705
1025 1705
0 3 34 0 0 8192 0 0 20 66 0 3
668 1698
668 1696
1025 1696
0 2 35 0 0 8192 0 0 20 61 0 3
516 1689
516 1687
1025 1687
0 4 33 0 0 8192 0 0 19 68 0 3
806 1647
806 1645
1024 1645
0 3 37 0 0 8192 0 0 19 94 0 3
699 1637
699 1636
1024 1636
0 2 35 0 0 0 0 0 19 61 0 3
516 1628
516 1627
1024 1627
0 4 36 0 0 0 0 0 18 92 0 3
844 1580
844 1579
1024 1579
0 3 37 0 0 0 0 0 18 94 0 2
699 1570
1024 1570
0 2 35 0 0 4096 0 0 18 82 0 3
516 2140
516 1561
1024 1561
0 4 33 0 0 0 0 0 17 68 0 2
806 1521
1022 1521
0 3 34 0 0 0 0 0 17 66 0 3
668 1513
668 1512
1022 1512
0 2 38 0 0 8192 0 0 17 96 0 3
547 1504
547 1503
1022 1503
0 4 36 0 0 0 0 0 16 92 0 2
844 1458
1020 1458
0 3 34 0 0 4224 0 0 16 87 0 3
668 2030
668 1449
1020 1449
0 2 38 0 0 0 0 0 16 96 0 3
547 1443
1020 1443
1020 1440
0 4 33 0 0 4224 0 0 15 89 0 3
806 1982
806 1394
1018 1394
0 3 37 0 0 0 0 0 15 94 0 3
699 1382
699 1385
1018 1385
0 2 38 0 0 0 0 0 15 96 0 4
547 1371
1014 1371
1014 1376
1018 1376
0 4 33 0 0 0 0 0 29 89 0 4
806 2341
996 2341
996 2326
1029 2326
0 3 34 0 0 0 0 0 29 87 0 4
668 2333
989 2333
989 2317
1029 2317
0 2 35 0 0 0 0 0 29 82 0 4
516 2324
982 2324
982 2308
1029 2308
0 4 36 0 0 0 0 0 28 93 0 4
844 2277
998 2277
998 2270
1028 2270
0 3 34 0 0 0 0 0 28 87 0 4
668 2268
992 2268
992 2261
1028 2261
0 2 35 0 0 0 0 0 28 82 0 4
516 2260
988 2260
988 2252
1028 2252
0 4 33 0 0 0 0 0 27 89 0 3
806 2217
1028 2217
1028 2214
0 3 37 0 0 8192 0 0 27 95 0 3
699 2207
699 2205
1028 2205
0 2 35 0 0 0 0 0 27 82 0 3
516 2198
516 2196
1028 2196
0 4 36 0 0 8192 0 0 26 93 0 3
844 2159
844 2158
1026 2158
0 3 37 0 0 0 0 0 26 95 0 2
699 2149
1026 2149
0 2 35 0 0 0 0 0 26 100 0 3
516 2451
516 2140
1026 2140
0 4 33 0 0 0 0 0 25 89 0 2
806 2101
1024 2101
0 3 34 0 0 0 0 0 25 87 0 3
668 2094
668 2092
1024 2092
0 2 38 0 0 8192 0 0 25 97 0 3
544 2084
544 2083
1024 2083
0 4 36 0 0 0 0 0 24 93 0 3
844 2041
844 2039
1024 2039
0 3 34 0 0 0 0 0 24 99 0 3
668 2441
668 2030
1024 2030
0 2 38 0 0 0 0 0 24 97 0 3
544 2022
544 2021
1024 2021
0 4 33 0 0 0 0 0 23 98 0 3
806 2436
806 1982
1024 1982
0 3 37 0 0 0 0 0 23 95 0 3
699 1974
699 1973
1024 1973
0 2 38 0 0 0 0 0 23 97 0 3
544 1963
544 1964
1024 1964
0 4 36 0 0 4224 0 0 14 93 0 3
844 1922
844 1327
1016 1327
2 4 36 0 0 0 0 32 22 0 0 3
844 2395
844 1922
1024 1922
0 3 37 0 0 4224 0 0 14 95 0 3
699 1914
699 1318
1016 1318
2 3 37 0 0 0 0 31 22 0 0 3
699 2400
699 1913
1024 1913
0 2 38 0 0 4224 0 0 14 97 0 3
547 1904
547 1309
1016 1309
2 2 38 0 0 0 0 30 22 0 0 3
544 2403
544 1904
1024 1904
1 1 33 0 0 0 0 5 32 0 0 3
790 2436
844 2436
844 2431
1 1 34 0 0 0 0 4 31 0 0 3
649 2441
699 2441
699 2436
1 1 35 0 0 0 0 3 30 0 0 3
502 2451
544 2451
544 2439
3 1 39 0 0 8320 0 40 39 0 0 3
1313 822
1385 822
1385 265
0 1 40 0 0 4224 0 0 55 103 0 3
926 1087
926 521
1014 521
1 1 40 0 0 0 0 66 47 0 0 5
1277 1148
1277 1163
923 1163
923 1087
1017 1087
1 0 2 0 0 0 0 48 0 0 105 3
1016 1031
904 1031
904 598
1 1 2 0 0 0 0 56 65 0 0 5
1013 466
904 466
904 598
1256 598
1256 602
2 1 41 0 0 8320 0 64 53 0 0 3
178 134
178 743
1012 743
0 1 4 0 0 0 0 0 64 110 0 3
134 135
134 134
142 134
2 1 42 0 0 4224 0 63 61 0 0 4
99 117
638 117
638 155
1006 155
0 1 5 0 0 0 0 0 63 111 0 3
62 89
63 89
63 117
1 1 4 0 0 0 0 7 54 0 0 3
134 37
134 683
1012 683
1 1 5 0 0 0 0 6 62 0 0 6
42 40
51 40
51 89
474 89
474 88
1004 88
5 1 43 0 0 4224 0 42 40 0 0 4
1189 806
1236 806
1236 813
1267 813
5 2 44 0 0 8320 0 41 40 0 0 4
1197 1002
1239 1002
1239 831
1267 831
0 0 45 0 0 8320 0 0 0 0 0 3
1275 880
1275 881
1272 881
5 4 46 0 0 4224 0 47 41 0 0 3
1062 1100
1147 1100
1147 1016
5 3 47 0 0 4224 0 48 41 0 0 4
1061 1044
1110 1044
1110 1007
1147 1007
5 2 48 0 0 12416 0 49 41 0 0 4
1061 988
1077 988
1077 998
1147 998
5 1 49 0 0 8320 0 50 41 0 0 4
1059 932
1108 932
1108 989
1147 989
5 4 50 0 0 8320 0 51 42 0 0 4
1057 875
1102 875
1102 820
1139 820
5 3 51 0 0 4224 0 52 42 0 0 4
1057 813
1122 813
1122 811
1139 811
5 2 52 0 0 12416 0 53 42 0 0 4
1057 756
1082 756
1082 802
1139 802
5 1 53 0 0 8320 0 54 42 0 0 4
1057 696
1095 696
1095 793
1139 793
3 1 54 0 0 4224 0 44 43 0 0 3
1255 272
1345 272
1345 266
5 2 55 0 0 8320 0 45 44 0 0 4
1178 402
1185 402
1185 281
1209 281
5 1 56 0 0 8320 0 46 44 0 0 4
1173 202
1190 202
1190 263
1209 263
5 4 57 0 0 8320 0 55 45 0 0 6
1059 534
1089 534
1089 439
1101 439
1101 416
1128 416
5 3 58 0 0 4224 0 56 45 0 0 5
1058 479
1058 426
1086 426
1086 407
1128 407
5 2 59 0 0 12416 0 57 45 0 0 4
1057 419
1076 419
1076 398
1128 398
0 1 60 0 0 4224 0 0 45 0 0 4
1060 354
1108 354
1108 389
1128 389
5 4 61 0 0 8320 0 59 46 0 0 4
1055 295
1082 295
1082 216
1123 216
5 3 62 0 0 12416 0 60 46 0 0 4
1053 232
1066 232
1066 207
1123 207
5 2 63 0 0 12416 0 61 46 0 0 4
1051 168
1082 168
1082 198
1123 198
5 1 64 0 0 8320 0 62 46 0 0 4
1049 101
1096 101
1096 189
1123 189
0 4 33 0 0 0 0 0 55 152 0 4
794 558
1007 558
1007 548
1014 548
0 3 34 0 0 0 0 0 55 150 0 4
656 548
1002 548
1002 539
1014 539
0 2 35 0 0 0 0 0 55 145 0 4
504 538
992 538
992 530
1014 530
0 4 36 0 0 0 0 0 56 176 0 3
832 494
832 493
1013 493
0 3 34 0 0 0 0 0 56 150 0 3
656 486
656 484
1013 484
0 2 35 0 0 0 0 0 56 145 0 3
504 477
504 475
1013 475
0 4 33 0 0 0 0 0 57 152 0 3
794 435
794 433
1012 433
0 3 37 0 0 0 0 0 57 178 0 3
687 425
687 424
1012 424
0 2 35 0 0 0 0 0 57 145 0 3
504 416
504 415
1012 415
0 4 36 0 0 0 0 0 58 176 0 3
832 368
832 367
1012 367
0 3 37 0 0 0 0 0 58 178 0 2
687 358
1012 358
0 2 35 0 0 0 0 0 58 166 0 3
504 928
504 349
1012 349
0 4 33 0 0 0 0 0 59 152 0 2
794 309
1010 309
0 3 34 0 0 0 0 0 59 150 0 3
656 301
656 300
1010 300
0 2 38 0 0 0 0 0 59 180 0 3
535 292
535 291
1010 291
0 4 36 0 0 0 0 0 60 176 0 2
832 246
1008 246
0 3 34 0 0 0 0 0 60 171 0 3
656 818
656 237
1008 237
0 2 38 0 0 0 0 0 60 180 0 3
535 231
1008 231
1008 228
0 4 33 0 0 0 0 0 61 173 0 3
794 770
794 182
1006 182
0 3 37 0 0 0 0 0 61 178 0 3
687 170
687 173
1006 173
0 2 38 0 0 0 0 0 61 180 0 4
535 159
1002 159
1002 164
1006 164
0 4 33 0 0 0 0 0 47 173 0 4
794 1129
984 1129
984 1114
1017 1114
0 3 34 0 0 0 0 0 47 171 0 4
656 1121
977 1121
977 1105
1017 1105
0 2 35 0 0 0 0 0 47 166 0 4
504 1112
970 1112
970 1096
1017 1096
0 4 36 0 0 0 0 0 48 177 0 4
832 1065
986 1065
986 1058
1016 1058
0 3 34 0 0 0 0 0 48 171 0 4
656 1056
980 1056
980 1049
1016 1049
0 2 35 0 0 0 0 0 48 166 0 4
504 1048
976 1048
976 1040
1016 1040
0 4 33 0 0 0 0 0 49 173 0 3
794 1005
1016 1005
1016 1002
0 3 37 0 0 0 0 0 49 179 0 3
687 995
687 993
1016 993
0 2 35 0 0 0 0 0 49 166 0 3
504 986
504 984
1016 984
0 4 36 0 0 0 0 0 50 177 0 3
832 947
832 946
1014 946
0 3 37 0 0 0 0 0 50 179 0 2
687 937
1014 937
0 2 35 0 0 8320 0 0 50 61 0 4
516 1561
504 1561
504 928
1014 928
0 4 33 0 0 0 0 0 51 173 0 2
794 889
1012 889
0 3 34 0 0 0 0 0 51 171 0 3
656 882
656 880
1012 880
0 2 38 0 0 0 0 0 51 181 0 3
532 872
532 871
1012 871
0 4 36 0 0 0 0 0 52 177 0 3
832 829
832 827
1012 827
0 3 34 0 0 0 0 0 52 66 0 5
671 1449
671 1229
656 1229
656 818
1012 818
0 2 38 0 0 0 0 0 52 181 0 3
532 810
532 809
1012 809
0 4 33 0 0 0 0 0 53 68 0 5
806 1397
806 1223
794 1223
794 770
1012 770
0 3 37 0 0 0 0 0 53 179 0 3
687 762
687 761
1012 761
0 2 38 0 0 0 0 0 53 181 0 3
532 751
532 752
1012 752
0 4 36 0 0 0 0 0 62 177 0 3
832 710
832 115
1004 115
0 4 36 0 0 0 0 0 54 92 0 5
844 1327
844 1183
832 1183
832 710
1012 710
0 3 37 0 0 0 0 0 62 179 0 3
687 702
687 106
1004 106
0 3 37 0 0 0 0 0 54 94 0 5
699 1320
699 1188
687 1188
687 701
1012 701
0 2 38 0 0 0 0 0 62 181 0 3
535 692
535 97
1004 97
0 2 38 0 0 0 0 0 54 96 0 5
547 1309
547 1284
532 1284
532 692
1012 692
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
