CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
71
13 Logic Switch~
5 230 2486 0 10 11
0 15 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43516 0
0
13 Logic Switch~
5 103 2489 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43516 1
0
13 Logic Switch~
5 244 1729 0 10 11
0 34 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43516 2
0
13 Logic Switch~
5 113 1733 0 10 11
0 35 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43516 3
0
13 Logic Switch~
5 200 883 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
43516 4
0
13 Logic Switch~
5 68 891 0 10 11
0 50 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
43516 5
0
13 Logic Switch~
5 143 214 0 10 11
0 64 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 B1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
43516 6
0
13 Logic Switch~
5 43 229 0 10 11
0 65 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7361 0 0
2
43516 7
0
13 Logic Switch~
5 356 46 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
43516 8
0
13 Logic Switch~
5 246 49 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
43516 9
0
13 Logic Switch~
5 137 54 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
43516 10
0
13 Logic Switch~
5 34 58 0 1 11
0 60
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
43516 11
0
14 Logic Display~
6 1019 83 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
43516 12
0
5 4071~
219 1017 3011 0 3 22
0 4 3 2
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U12D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 12 0
1 U
4597 0 0
2
43516 13
0
5 4081~
219 896 3070 0 3 22
0 6 5 3
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U14D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 14 0
1 U
3835 0 0
2
43516 14
0
5 4081~
219 892 2967 0 3 22
0 8 7 4
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U14C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 14 0
1 U
3670 0 0
2
43516 15
0
14 Logic Display~
6 1146 83 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
43516 16
0
5 4030~
219 994 2722 0 3 22
0 8 7 9
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U11D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 11 0
1 U
9323 0 0
2
43516 17
0
5 4030~
219 867 2613 0 3 22
0 6 5 8
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U11C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
317 0 0
2
43516 18
0
5 4081~
219 601 2866 0 3 22
0 11 10 7
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U14B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 14 0
1 U
3108 0 0
2
43516 19
0
5 4049~
219 307 2768 0 2 22
0 15 14
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
4299 0 0
2
43516 20
0
5 4071~
219 678 2711 0 3 22
0 13 12 5
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U12C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 12 0
1 U
9672 0 0
2
43516 21
0
5 4081~
219 598 2754 0 3 22
0 16 14 12
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U14A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 14 0
1 U
7876 0 0
2
43516 22
0
5 4081~
219 598 2682 0 3 22
0 17 15 13
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 10 0
1 U
6369 0 0
2
43516 23
0
5 4071~
219 678 2584 0 3 22
0 19 18 6
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 12 0
1 U
9172 0 0
2
43516 24
0
5 4073~
219 599 2540 0 4 22
0 20 21 22 19
0
0 0 624 0
4 4073
-7 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 13 0
1 U
7100 0 0
2
43516 25
0
5 4030~
219 428 2512 0 3 22
0 16 15 22
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U11B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
3820 0 0
2
43516 26
0
5 4071~
219 1104 2312 0 3 22
0 24 23 10
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U12A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 12 0
1 U
7678 0 0
2
43516 27
0
5 4081~
219 1001 2368 0 3 22
0 26 25 23
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 10 0
1 U
961 0 0
2
43516 28
0
5 4081~
219 996 2286 0 3 22
0 28 27 24
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
3178 0 0
2
43516 29
0
14 Logic Display~
6 1191 87 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
43516 30
0
5 4030~
219 982 1954 0 3 22
0 28 27 29
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U11A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
3951 0 0
2
43516 31
0
5 4030~
219 869 1881 0 3 22
0 26 25 28
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U8D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
8885 0 0
2
43516 32
0
5 4049~
219 356 2049 0 2 22
0 34 33
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
3780 0 0
2
43516 33
0
5 4081~
219 596 2206 0 3 22
0 30 11 27
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U10A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
9265 0 0
2
43516 34
0
5 4071~
219 688 1998 0 3 22
0 32 31 25
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
9442 0 0
2
43516 35
0
5 4081~
219 598 2046 0 3 22
0 16 33 31
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 9 0
1 U
9424 0 0
2
43516 36
0
5 4081~
219 599 1962 0 3 22
0 17 34 32
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
9968 0 0
2
43516 37
0
5 4071~
219 682 1841 0 3 22
0 36 35 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
9281 0 0
2
43516 38
0
5 4073~
219 602 1792 0 4 22
0 20 21 37 36
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
8464 0 0
2
43516 39
0
5 4030~
219 472 1761 0 3 22
0 16 34 37
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U8C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
7168 0 0
2
43516 40
0
5 4071~
219 998 1454 0 3 22
0 39 38 30
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
3171 0 0
2
43516 41
0
5 4081~
219 917 1509 0 3 22
0 41 40 38
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
4139 0 0
2
43516 42
0
5 4081~
219 913 1417 0 3 22
0 43 42 39
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U9A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
6435 0 0
2
43516 43
0
14 Logic Display~
6 1233 89 0 1 2
10 44
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
43516 44
0
5 4030~
219 967 1126 0 3 22
0 43 42 44
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U8B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
6874 0 0
2
43516 45
0
5 4030~
219 887 1012 0 3 22
0 41 40 43
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U8A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 8 0
1 U
5305 0 0
2
43516 46
0
5 4081~
219 624 1320 0 3 22
0 11 45 42
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
34 0 0
2
43516 47
0
5 4049~
219 230 1000 0 2 22
0 49 48
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
969 0 0
2
43516 48
0
5 4071~
219 713 1138 0 3 22
0 47 46 40
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
8402 0 0
2
43516 49
0
5 4081~
219 626 1196 0 3 22
0 16 48 46
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
3751 0 0
2
43516 50
0
5 4081~
219 628 1099 0 3 22
0 17 49 47
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
4292 0 0
2
43516 51
0
5 4071~
219 713 961 0 3 22
0 51 50 41
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
6118 0 0
2
43516 52
0
5 4073~
219 630 919 0 4 22
0 20 21 52 51
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 2 0
1 U
34 0 0
2
43516 53
0
5 4030~
219 492 901 0 3 22
0 16 49 52
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
6357 0 0
2
43516 54
0
5 4071~
219 1094 610 0 3 22
0 54 53 45
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
319 0 0
2
43516 55
0
5 4081~
219 1023 656 0 3 22
0 56 55 53
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
3976 0 0
2
43516 56
0
5 4081~
219 1023 581 0 3 22
0 57 58 54
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
7634 0 0
2
43516 57
0
5 4030~
219 1047 308 0 3 22
0 57 58 59
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
523 0 0
2
43516 58
0
14 Logic Display~
6 1282 91 0 1 2
10 59
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
43516 59
0
5 4030~
219 917 248 0 3 22
0 56 55 57
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
6901 0 0
2
43516 60
0
5 4049~
219 204 167 0 2 22
0 21 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
842 0 0
2
43516 61
0
5 4081~
219 722 488 0 3 22
0 11 60 58
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
3277 0 0
2
43516 62
0
5 4049~
219 218 367 0 2 22
0 64 63
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
4212 0 0
2
43516 63
0
5 4081~
219 724 392 0 3 22
0 16 63 61
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
4720 0 0
2
43516 64
0
5 4071~
219 812 360 0 3 22
0 62 61 55
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
5551 0 0
2
43516 65
0
5 4081~
219 721 329 0 3 22
0 17 64 62
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
6986 0 0
2
43516 66
0
5 4071~
219 803 210 0 3 22
0 66 65 56
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
8745 0 0
2
43516 67
0
5 4049~
219 420 70 0 2 22
0 17 20
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U3A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
9592 0 0
2
43516 68
0
5 4073~
219 721 189 0 4 22
0 67 21 20 66
0
0 0 624 0
4 4073
-7 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
8748 0 0
2
43516 69
0
5 4030~
219 557 180 0 3 22
0 16 64 67
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
7168 0 0
2
43516 70
0
111
3 1 2 0 0 8320 0 14 13 0 0 5
1050 3011
1312 3011
1312 142
1019 142
1019 101
3 2 3 0 0 4224 0 15 14 0 0 4
917 3070
972 3070
972 3020
1004 3020
3 1 4 0 0 12416 0 16 14 0 0 4
913 2967
952 2967
952 3002
1004 3002
0 2 5 0 0 4224 0 0 15 11 0 3
718 2711
718 3079
872 3079
0 1 6 0 0 4224 0 0 15 12 0 3
759 2584
759 3061
872 3061
0 2 7 0 0 8192 0 0 16 9 0 3
736 2866
736 2976
868 2976
0 1 8 0 0 8320 0 0 16 10 0 4
920 2712
857 2712
857 2958
868 2958
1 3 9 0 0 4224 0 17 18 0 0 3
1146 101
1146 2722
1027 2722
3 2 7 0 0 4224 0 20 18 0 0 4
622 2866
834 2866
834 2731
978 2731
3 1 8 0 0 0 0 19 18 0 0 4
900 2613
920 2613
920 2713
978 2713
3 2 5 0 0 0 0 22 19 0 0 4
711 2711
819 2711
819 2622
851 2622
3 1 6 0 0 0 0 25 19 0 0 4
711 2584
812 2584
812 2604
851 2604
3 2 10 0 0 12416 0 28 20 0 0 10
1137 2312
1150 2312
1150 2447
793 2447
793 2803
497 2803
497 2878
554 2878
554 2875
577 2875
0 1 11 0 0 4096 0 0 20 40 0 3
342 2215
342 2857
577 2857
3 2 12 0 0 12416 0 23 22 0 0 4
619 2754
629 2754
629 2720
665 2720
3 1 13 0 0 4224 0 24 22 0 0 4
619 2682
649 2682
649 2702
665 2702
2 2 14 0 0 4224 0 21 23 0 0 4
328 2768
559 2768
559 2763
574 2763
0 1 15 0 0 8192 0 0 21 21 0 4
292 2691
259 2691
259 2768
292 2768
0 1 16 0 0 4096 0 0 23 27 0 3
332 2503
332 2745
574 2745
0 1 17 0 0 4096 0 0 24 47 0 5
437 1953
437 2421
556 2421
556 2673
574 2673
0 2 15 0 0 8320 0 0 24 28 0 3
292 2521
292 2691
574 2691
1 2 18 0 0 12416 0 2 25 0 0 6
115 2489
130 2489
130 2596
613 2596
613 2593
665 2593
4 1 19 0 0 8320 0 26 25 0 0 4
620 2540
643 2540
643 2575
665 2575
0 1 20 0 0 8192 0 0 26 51 0 6
451 1687
418 1687
418 2457
500 2457
500 2531
575 2531
0 2 21 0 0 12288 0 0 26 52 0 7
356 1707
356 1964
389 1964
389 2471
490 2471
490 2540
575 2540
3 3 22 0 0 12416 0 27 26 0 0 4
461 2512
479 2512
479 2549
575 2549
0 1 16 0 0 4096 0 0 27 44 0 5
282 2013
282 2466
311 2466
311 2503
412 2503
1 2 15 0 0 0 0 1 27 0 0 4
242 2486
282 2486
282 2521
412 2521
3 2 23 0 0 8320 0 29 28 0 0 4
1022 2368
1049 2368
1049 2321
1091 2321
3 1 24 0 0 12416 0 30 28 0 0 4
1017 2286
1044 2286
1044 2303
1091 2303
0 2 25 0 0 4224 0 0 29 38 0 3
738 1998
738 2377
977 2377
0 1 26 0 0 4224 0 0 29 39 0 3
773 1841
773 2359
977 2359
0 2 27 0 0 8192 0 0 30 36 0 3
807 2206
807 2295
972 2295
0 1 28 0 0 4224 0 0 30 37 0 3
923 1945
923 2277
972 2277
1 3 29 0 0 4224 0 31 32 0 0 3
1191 105
1191 1954
1015 1954
3 2 27 0 0 4224 0 35 32 0 0 4
617 2206
906 2206
906 1963
966 1963
3 1 28 0 0 0 0 33 32 0 0 4
902 1881
914 1881
914 1945
966 1945
3 2 25 0 0 0 0 36 33 0 0 4
721 1998
747 1998
747 1890
853 1890
3 1 26 0 0 0 0 39 33 0 0 4
715 1841
828 1841
828 1872
853 1872
0 2 11 0 0 4096 0 0 35 68 0 3
306 1311
306 2215
572 2215
3 1 30 0 0 16512 0 42 35 0 0 8
1031 1454
1072 1454
1072 1589
811 1589
811 2153
496 2153
496 2197
572 2197
3 2 31 0 0 8320 0 37 36 0 0 4
619 2046
639 2046
639 2007
675 2007
3 1 32 0 0 12416 0 38 36 0 0 4
620 1962
634 1962
634 1989
675 1989
0 1 16 0 0 0 0 0 37 55 0 5
282 1664
282 2013
514 2013
514 2037
574 2037
2 2 33 0 0 4224 0 34 37 0 0 4
377 2049
511 2049
511 2055
574 2055
0 1 34 0 0 4096 0 0 34 48 0 3
330 1971
330 2049
341 2049
0 1 17 0 0 4224 0 0 38 75 0 3
383 1090
383 1953
575 1953
0 2 34 0 0 8320 0 0 38 54 0 3
313 1770
313 1971
575 1971
1 2 35 0 0 12416 0 4 39 0 0 4
125 1733
166 1733
166 1850
669 1850
4 1 36 0 0 8320 0 40 39 0 0 4
623 1792
641 1792
641 1832
669 1832
0 1 20 0 0 4224 0 0 40 78 0 5
451 847
451 1694
553 1694
553 1783
578 1783
0 2 21 0 0 4224 0 0 40 79 0 5
356 863
356 1707
526 1707
526 1792
578 1792
3 3 37 0 0 12416 0 41 40 0 0 4
505 1761
516 1761
516 1801
578 1801
1 2 34 0 0 0 0 3 41 0 0 4
256 1729
313 1729
313 1770
456 1770
0 1 16 0 0 4096 0 0 41 73 0 5
267 1187
267 1664
361 1664
361 1752
456 1752
3 2 38 0 0 8320 0 43 42 0 0 4
938 1509
958 1509
958 1463
985 1463
3 1 39 0 0 12416 0 44 42 0 0 4
934 1417
951 1417
951 1445
985 1445
0 2 40 0 0 4224 0 0 43 65 0 3
752 1138
752 1518
893 1518
0 1 41 0 0 4224 0 0 43 66 0 3
764 961
764 1500
893 1500
0 2 42 0 0 8192 0 0 44 64 0 3
776 1320
776 1426
889 1426
0 1 43 0 0 4224 0 0 44 63 0 5
920 1117
920 1337
860 1337
860 1408
889 1408
1 3 44 0 0 4224 0 45 46 0 0 3
1233 107
1233 1126
1000 1126
3 1 43 0 0 0 0 47 46 0 0 3
920 1012
920 1117
951 1117
3 2 42 0 0 4224 0 48 46 0 0 4
645 1320
837 1320
837 1135
951 1135
3 2 40 0 0 0 0 50 47 0 0 4
746 1138
811 1138
811 1021
871 1021
3 1 41 0 0 0 0 53 47 0 0 4
746 961
829 961
829 1003
871 1003
3 2 45 0 0 16512 0 56 48 0 0 8
1127 610
1140 610
1140 778
781 778
781 1274
526 1274
526 1329
600 1329
0 1 11 0 0 4224 0 0 48 95 0 3
291 318
291 1311
600 1311
3 2 46 0 0 8320 0 51 50 0 0 4
647 1196
686 1196
686 1147
700 1147
3 1 47 0 0 4224 0 52 50 0 0 4
649 1099
681 1099
681 1129
700 1129
2 2 48 0 0 12416 0 49 51 0 0 4
251 1000
256 1000
256 1205
602 1205
0 1 49 0 0 8192 0 0 49 81 0 4
212 909
200 909
200 1000
215 1000
0 1 16 0 0 0 0 0 51 82 0 3
267 892
267 1187
602 1187
0 2 49 0 0 8320 0 0 52 81 0 3
324 910
324 1108
604 1108
0 1 17 0 0 0 0 0 52 103 0 3
383 320
383 1090
604 1090
1 2 50 0 0 12416 0 6 53 0 0 4
80 891
112 891
112 970
700 970
4 1 51 0 0 8320 0 54 53 0 0 4
651 919
680 919
680 952
700 952
0 1 20 0 0 0 0 0 54 106 0 5
451 70
451 847
594 847
594 910
606 910
0 2 21 0 0 0 0 0 54 108 0 5
356 231
356 863
580 863
580 919
606 919
3 3 52 0 0 12416 0 55 54 0 0 4
525 901
550 901
550 928
606 928
1 2 49 0 0 0 0 5 55 0 0 3
212 883
212 910
476 910
0 1 16 0 0 4224 0 0 55 101 0 3
267 383
267 892
476 892
3 2 53 0 0 8320 0 57 56 0 0 4
1044 656
1051 656
1051 619
1081 619
3 1 54 0 0 4224 0 58 56 0 0 4
1044 581
1066 581
1066 601
1081 601
0 2 55 0 0 4224 0 0 57 92 0 3
871 360
871 665
999 665
0 1 56 0 0 4224 0 0 57 93 0 3
858 210
858 647
999 647
0 1 57 0 0 4224 0 0 58 91 0 3
963 248
963 572
999 572
0 2 58 0 0 8320 0 0 58 90 0 3
803 488
803 590
999 590
3 1 59 0 0 4224 0 59 60 0 0 3
1080 308
1282 308
1282 109
3 2 58 0 0 0 0 63 59 0 0 4
743 488
923 488
923 317
1031 317
3 1 57 0 0 0 0 61 59 0 0 4
950 248
988 248
988 299
1031 299
3 2 55 0 0 0 0 66 61 0 0 4
845 360
877 360
877 257
901 257
3 1 56 0 0 0 0 68 61 0 0 4
836 210
884 210
884 239
901 239
1 2 60 0 0 12416 0 12 63 0 0 4
46 58
76 58
76 497
698 497
2 1 11 0 0 0 0 62 63 0 0 5
225 167
225 318
330 318
330 479
698 479
0 1 21 0 0 0 0 0 62 108 0 3
171 140
171 167
189 167
3 2 61 0 0 12416 0 65 66 0 0 4
745 392
766 392
766 369
799 369
3 1 62 0 0 12416 0 67 66 0 0 4
742 329
764 329
764 351
799 351
2 2 63 0 0 12416 0 64 65 0 0 4
239 367
258 367
258 401
700 401
0 1 64 0 0 4096 0 0 64 102 0 3
179 338
179 367
203 367
0 1 16 0 0 0 0 0 65 111 0 3
267 171
267 383
700 383
0 2 64 0 0 8320 0 0 67 110 0 3
179 214
179 338
697 338
0 1 17 0 0 0 0 0 67 107 0 3
383 46
383 320
697 320
1 2 65 0 0 12416 0 8 68 0 0 6
55 229
91 229
91 256
759 256
759 219
790 219
4 1 66 0 0 4224 0 70 68 0 0 4
742 189
779 189
779 201
790 201
2 3 20 0 0 0 0 69 70 0 0 4
441 70
621 70
621 198
697 198
1 1 17 0 0 0 0 9 69 0 0 4
368 46
398 46
398 70
405 70
1 2 21 0 0 0 0 11 70 0 0 7
149 54
149 140
251 140
251 231
592 231
592 189
697 189
3 1 67 0 0 4224 0 71 70 0 0 2
590 180
697 180
1 2 64 0 0 0 0 7 71 0 0 4
155 214
409 214
409 189
541 189
1 1 16 0 0 0 0 10 71 0 0 4
258 49
267 49
267 171
541 171
2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 5
1000 26 1036 42
1000 26 1036 42
5 Carry
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 32768 0 2
1259 32 1275 48
1259 32 1275 48
2 F1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
