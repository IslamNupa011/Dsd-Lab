CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 506 1251 0 10 11
0 33 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9424 0 0
2
5.89879e-315 5.41378e-315
0
13 Logic Switch~
5 653 1241 0 1 11
0 32
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 s1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9968 0 0
2
5.89879e-315 5.4086e-315
0
13 Logic Switch~
5 794 1236 0 1 11
0 31
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9281 0 0
2
5.89879e-315 5.40342e-315
0
13 Logic Switch~
5 150 49 0 10 11
0 7 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8464 0 0
2
5.89879e-315 0
0
13 Logic Switch~
5 58 52 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 A0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7168 0 0
2
5.89879e-315 0
0
14 Logic Display~
6 1408 261 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3171 0 0
2
43493 0
0
2 +V
167 1305 1151 0 1 3
0 5
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89879e-315 0
0
7 Ground~
168 1284 620 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
5.89879e-315 0
0
5 4049~
219 185 146 0 2 22
0 7 8
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 9 0
1 U
5283 0 0
2
5.89879e-315 0
0
5 4049~
219 106 129 0 2 22
0 6 9
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 9 0
1 U
6874 0 0
2
5.89879e-315 0
0
5 4082~
219 1056 113 0 5 22
0 6 36 35 34 30
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
5305 0 0
2
5.89879e-315 5.463e-315
0
5 4082~
219 1058 180 0 5 22
0 9 36 35 31 29
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U1B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 1 0
1 U
34 0 0
2
5.89879e-315 5.46041e-315
0
5 4082~
219 1060 244 0 5 22
0 2 36 32 34 28
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
969 0 0
2
5.89879e-315 5.45782e-315
0
5 4082~
219 1062 307 0 5 22
0 7 36 32 31 27
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U2B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
8402 0 0
2
5.89879e-315 5.45523e-315
0
5 4082~
219 1064 365 0 5 22
0 7 33 35 34 4
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
3751 0 0
2
5.89879e-315 5.45264e-315
0
5 4082~
219 1064 431 0 5 22
0 7 33 35 31 26
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
4292 0 0
2
5.89879e-315 5.45005e-315
0
5 4082~
219 1065 491 0 5 22
0 2 33 32 34 25
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
6118 0 0
2
5.89879e-315 5.44746e-315
0
5 4082~
219 1066 546 0 5 22
0 5 33 32 31 24
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U4B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
34 0 0
2
5.89879e-315 5.44487e-315
0
5 4082~
219 1064 708 0 5 22
0 7 36 35 34 20
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
6357 0 0
2
5.89879e-315 5.44228e-315
0
5 4082~
219 1064 768 0 5 22
0 8 36 35 31 19
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U5B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
319 0 0
2
5.89879e-315 5.43969e-315
0
5 4082~
219 1064 825 0 5 22
0 6 36 32 34 18
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 6 0
1 U
3976 0 0
2
5.89879e-315 5.4371e-315
0
5 4082~
219 1064 887 0 5 22
0 2 36 32 31 17
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U6B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 6 0
1 U
7634 0 0
2
5.89879e-315 5.43451e-315
0
5 4082~
219 1066 944 0 5 22
0 6 33 35 34 16
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 7 0
1 U
523 0 0
2
5.89879e-315 5.43192e-315
0
5 4082~
219 1068 1000 0 5 22
0 6 33 35 31 15
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U7B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 7 0
1 U
6748 0 0
2
5.89879e-315 5.42933e-315
0
5 4082~
219 1068 1056 0 5 22
0 2 33 32 34 14
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
6901 0 0
2
5.89879e-315 5.42414e-315
0
5 4082~
219 1069 1112 0 5 22
0 5 33 32 31 13
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U8B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
842 0 0
2
5.89879e-315 5.41896e-315
0
5 4049~
219 557 1221 0 2 22
0 33 36
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9A
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 9 0
1 U
3277 0 0
2
5.89879e-315 5.39824e-315
0
5 4049~
219 712 1218 0 2 22
0 32 35
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9B
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 9 0
1 U
4212 0 0
2
5.89879e-315 5.39306e-315
0
5 4049~
219 857 1213 0 2 22
0 31 34
0
0 0 624 90
4 4049
-7 -24 21 -16
3 U9C
16 -2 37 6
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 9 0
1 U
4720 0 0
2
5.89879e-315 5.38788e-315
0
8 4-In OR~
219 1168 214 0 5 22
0 30 29 28 27 23
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 10 0
1 U
5551 0 0
2
5.89879e-315 5.37752e-315
0
8 4-In OR~
219 1173 414 0 5 22
0 4 26 25 24 22
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U10B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 10 0
1 U
6986 0 0
2
5.89879e-315 5.36716e-315
0
5 4071~
219 1250 284 0 3 22
0 23 22 21
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
8745 0 0
2
5.89879e-315 5.3568e-315
0
14 Logic Display~
6 1373 260 0 1 2
10 21
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9592 0 0
2
5.89879e-315 5.34643e-315
0
8 4-In OR~
219 1184 818 0 5 22
0 20 19 18 17 10
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 12 0
1 U
8748 0 0
2
5.89879e-315 5.32571e-315
0
8 4-In OR~
219 1192 1014 0 5 22
0 16 15 14 13 11
0
0 0 624 0
4 4072
-14 -24 14 -16
4 U12B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 12 0
1 U
7168 0 0
2
5.89879e-315 5.30499e-315
0
5 4071~
219 1308 834 0 3 22
0 10 11 3
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
631 0 0
2
5.89879e-315 5.26354e-315
0
92
3 1 3 0 0 8320 0 36 6 0 0 3
1341 834
1408 834
1408 279
1 5 4 0 0 4224 0 31 15 0 0 4
1156 401
1115 401
1115 365
1085 365
0 1 5 0 0 4224 0 0 18 4 0 3
954 1099
954 533
1042 533
1 1 5 0 0 0 0 7 26 0 0 5
1305 1160
1305 1175
951 1175
951 1099
1045 1099
1 0 2 0 0 8192 0 25 0 0 6 3
1044 1043
932 1043
932 610
1 0 2 0 0 0 0 17 0 0 13 3
1041 478
932 478
932 610
1 0 6 0 0 4224 0 24 0 0 9 3
1044 987
80 987
80 931
1 0 7 0 0 4224 0 16 0 0 19 2
1040 418
162 418
1 0 6 0 0 0 0 23 0 0 14 3
1042 931
79 931
79 807
1 0 7 0 0 0 0 15 0 0 19 2
1040 352
162 352
1 0 2 0 0 4096 0 22 0 0 13 3
1040 874
140 874
140 610
1 0 7 0 0 0 0 14 0 0 19 2
1038 294
162 294
1 1 2 0 0 8320 0 8 13 0 0 5
1284 614
1284 610
132 610
132 231
1036 231
0 1 6 0 0 0 0 0 21 20 0 3
79 100
79 812
1040 812
2 1 8 0 0 8320 0 9 20 0 0 3
206 146
206 755
1040 755
0 1 7 0 0 0 0 0 9 19 0 3
162 147
162 146
170 146
2 1 9 0 0 4224 0 10 12 0 0 4
127 129
666 129
666 167
1034 167
0 1 6 0 0 0 0 0 10 20 0 3
90 101
91 101
91 129
1 1 7 0 0 0 0 4 19 0 0 3
162 49
162 695
1040 695
1 1 6 0 0 0 0 5 11 0 0 6
70 52
79 52
79 101
502 101
502 100
1032 100
5 1 10 0 0 4224 0 34 36 0 0 4
1217 818
1264 818
1264 825
1295 825
5 2 11 0 0 8320 0 35 36 0 0 4
1225 1014
1267 1014
1267 843
1295 843
0 0 12 0 0 8320 0 0 0 0 0 3
1303 892
1303 893
1300 893
5 4 13 0 0 4224 0 26 35 0 0 3
1090 1112
1175 1112
1175 1028
5 3 14 0 0 4224 0 25 35 0 0 4
1089 1056
1138 1056
1138 1019
1175 1019
5 2 15 0 0 12416 0 24 35 0 0 4
1089 1000
1105 1000
1105 1010
1175 1010
5 1 16 0 0 8320 0 23 35 0 0 4
1087 944
1136 944
1136 1001
1175 1001
5 4 17 0 0 8320 0 22 34 0 0 4
1085 887
1130 887
1130 832
1167 832
5 3 18 0 0 4224 0 21 34 0 0 4
1085 825
1150 825
1150 823
1167 823
5 2 19 0 0 12416 0 20 34 0 0 4
1085 768
1110 768
1110 814
1167 814
5 1 20 0 0 8320 0 19 34 0 0 4
1085 708
1123 708
1123 805
1167 805
3 1 21 0 0 4224 0 32 33 0 0 3
1283 284
1373 284
1373 278
5 2 22 0 0 8320 0 31 32 0 0 4
1206 414
1213 414
1213 293
1237 293
5 1 23 0 0 8320 0 30 32 0 0 4
1201 214
1218 214
1218 275
1237 275
5 4 24 0 0 8320 0 18 31 0 0 6
1087 546
1117 546
1117 451
1129 451
1129 428
1156 428
5 3 25 0 0 4224 0 17 31 0 0 5
1086 491
1086 438
1114 438
1114 419
1156 419
5 2 26 0 0 12416 0 16 31 0 0 4
1085 431
1104 431
1104 410
1156 410
5 4 27 0 0 8320 0 14 30 0 0 4
1083 307
1110 307
1110 228
1151 228
5 3 28 0 0 12416 0 13 30 0 0 4
1081 244
1094 244
1094 219
1151 219
5 2 29 0 0 12416 0 12 30 0 0 4
1079 180
1110 180
1110 210
1151 210
5 1 30 0 0 8320 0 11 30 0 0 4
1077 113
1124 113
1124 201
1151 201
0 4 31 0 0 4096 0 0 18 60 0 4
822 570
1035 570
1035 560
1042 560
0 3 32 0 0 4096 0 0 18 58 0 4
684 560
1030 560
1030 551
1042 551
0 2 33 0 0 4096 0 0 18 53 0 4
532 550
1020 550
1020 542
1042 542
0 4 34 0 0 8192 0 0 17 84 0 3
860 506
860 505
1041 505
0 3 32 0 0 8192 0 0 17 58 0 3
684 498
684 496
1041 496
0 2 33 0 0 8192 0 0 17 53 0 3
532 489
532 487
1041 487
0 4 31 0 0 8192 0 0 16 60 0 3
822 447
822 445
1040 445
0 3 35 0 0 8192 0 0 16 86 0 3
715 437
715 436
1040 436
0 2 33 0 0 0 0 0 16 53 0 3
532 428
532 427
1040 427
0 4 34 0 0 0 0 0 15 84 0 3
860 380
860 379
1040 379
0 3 35 0 0 0 0 0 15 86 0 2
715 370
1040 370
0 2 33 0 0 4224 0 0 15 74 0 3
532 940
532 361
1040 361
0 4 31 0 0 0 0 0 14 60 0 2
822 321
1038 321
0 3 32 0 0 0 0 0 14 58 0 3
684 313
684 312
1038 312
0 2 36 0 0 8192 0 0 14 88 0 3
563 304
563 303
1038 303
0 4 34 0 0 0 0 0 13 84 0 2
860 258
1036 258
0 3 32 0 0 4224 0 0 13 79 0 3
684 830
684 249
1036 249
0 2 36 0 0 0 0 0 13 88 0 3
563 243
1036 243
1036 240
0 4 31 0 0 4224 0 0 12 81 0 3
822 782
822 194
1034 194
0 3 35 0 0 0 0 0 12 86 0 3
715 182
715 185
1034 185
0 2 36 0 0 0 0 0 12 88 0 4
563 171
1030 171
1030 176
1034 176
0 4 31 0 0 0 0 0 26 81 0 4
822 1141
1012 1141
1012 1126
1045 1126
0 3 32 0 0 0 0 0 26 79 0 4
684 1133
1005 1133
1005 1117
1045 1117
0 2 33 0 0 0 0 0 26 74 0 4
532 1124
998 1124
998 1108
1045 1108
0 4 34 0 0 0 0 0 25 85 0 4
860 1077
1014 1077
1014 1070
1044 1070
0 3 32 0 0 0 0 0 25 79 0 4
684 1068
1008 1068
1008 1061
1044 1061
0 2 33 0 0 0 0 0 25 74 0 4
532 1060
1004 1060
1004 1052
1044 1052
0 4 31 0 0 0 0 0 24 81 0 3
822 1017
1044 1017
1044 1014
0 3 35 0 0 8192 0 0 24 87 0 3
715 1007
715 1005
1044 1005
0 2 33 0 0 0 0 0 24 74 0 3
532 998
532 996
1044 996
0 4 34 0 0 8192 0 0 23 85 0 3
860 959
860 958
1042 958
0 3 35 0 0 0 0 0 23 87 0 2
715 949
1042 949
0 2 33 0 0 0 0 0 23 92 0 3
532 1251
532 940
1042 940
0 4 31 0 0 0 0 0 22 81 0 2
822 901
1040 901
0 3 32 0 0 0 0 0 22 79 0 3
684 894
684 892
1040 892
0 2 36 0 0 8192 0 0 22 89 0 3
560 884
560 883
1040 883
0 4 34 0 0 0 0 0 21 85 0 3
860 841
860 839
1040 839
0 3 32 0 0 0 0 0 21 91 0 3
684 1241
684 830
1040 830
0 2 36 0 0 0 0 0 21 89 0 3
560 822
560 821
1040 821
0 4 31 0 0 0 0 0 20 90 0 3
822 1236
822 782
1040 782
0 3 35 0 0 0 0 0 20 87 0 3
715 774
715 773
1040 773
0 2 36 0 0 0 0 0 20 89 0 3
560 763
560 764
1040 764
0 4 34 0 0 4224 0 0 11 85 0 3
860 722
860 127
1032 127
2 4 34 0 0 0 0 29 19 0 0 3
860 1195
860 722
1040 722
0 3 35 0 0 4224 0 0 11 87 0 3
715 714
715 118
1032 118
2 3 35 0 0 0 0 28 19 0 0 3
715 1200
715 713
1040 713
0 2 36 0 0 4224 0 0 11 89 0 3
563 704
563 109
1032 109
2 2 36 0 0 0 0 27 19 0 0 3
560 1203
560 704
1040 704
1 1 31 0 0 0 0 3 29 0 0 3
806 1236
860 1236
860 1231
1 1 32 0 0 0 0 2 28 0 0 3
665 1241
715 1241
715 1236
1 1 33 0 0 0 0 1 27 0 0 3
518 1251
560 1251
560 1239
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
