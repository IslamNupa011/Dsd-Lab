CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 699 79 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 CPi
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5283 0 0
2
43550.5 0
0
13 Logic Switch~
5 913 286 0 10 11
0 24 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 reset
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6874 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 91 72 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 P5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5305 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 195 73 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
34 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 280 81 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
969 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 362 84 0 1 11
0 16
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8402 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 435 88 0 1 11
0 5
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 P1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3751 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 499 93 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
1 B
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4292 0 0
2
5.89886e-315 0
0
13 Logic Switch~
5 564 99 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -15 9 -7
1 C
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6118 0 0
2
5.89886e-315 0
0
14 Logic Display~
6 999 80 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
34 0 0
2
43550.5 0
0
5 4081~
219 881 630 0 3 22
0 6 5 4
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
6357 0 0
2
43550.5 0
0
5 4071~
219 798 614 0 3 22
0 8 7 6
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
319 0 0
2
43550.5 0
0
5 4081~
219 729 645 0 3 22
0 10 9 7
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
3976 0 0
2
43550.5 0
0
5 4081~
219 728 586 0 3 22
0 12 11 8
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
7634 0 0
2
43550.5 0
0
5 4030~
219 646 566 0 3 22
0 10 9 12
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U2B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
523 0 0
2
43550.5 0
0
8 4-In OR~
219 735 462 0 5 22
0 17 14 16 15 13
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5B
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 5 0
1 U
6748 0 0
2
43550.5 0
0
5 4081~
219 657 458 0 3 22
0 9 18 14
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
6901 0 0
2
43550.5 0
0
8 4-In OR~
219 716 335 0 5 22
0 17 21 20 18 19
0
0 0 624 0
4 4072
-14 -24 14 -16
3 U5A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 5 0
1 U
842 0 0
2
43550.5 0
0
5 4081~
219 585 359 0 3 22
0 22 15 21
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
3277 0 0
2
43550.5 0
0
5 4049~
219 521 334 0 2 22
0 9 22
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 4 0
1 U
4212 0 0
2
43550.5 0
0
5 4081~
219 628 279 0 3 22
0 23 5 17
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
4720 0 0
2
43550.5 0
0
5 4030~
219 560 228 0 3 22
0 9 11 23
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U2A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
5551 0 0
2
43550.5 0
0
14 Logic Display~
6 1114 80 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6986 0 0
2
5.89886e-315 0
0
7 Pulser~
4 778 202 0 11 12
0 3 25 2 26 0 0 5 5 -1
7 1
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8745 0 0
2
5.89886e-315 0
0
6 JK RN~
219 919 193 0 6 22
0 19 2 13 24 27 10
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9592 0 0
2
5.89886e-315 0
0
34
3 2 2 0 0 12416 0 24 25 0 0 4
802 193
822 193
822 185
888 185
1 1 3 0 0 4224 0 1 24 0 0 3
711 79
711 193
754 193
1 3 4 0 0 4224 0 10 11 0 0 3
999 98
999 630
902 630
0 2 5 0 0 8320 0 0 11 29 0 5
447 288
447 672
835 672
835 639
857 639
3 1 6 0 0 12416 0 12 11 0 0 4
831 614
837 614
837 621
857 621
3 2 7 0 0 8320 0 13 12 0 0 4
750 645
765 645
765 623
785 623
3 1 8 0 0 8320 0 14 12 0 0 3
749 586
749 605
785 605
0 2 9 0 0 8192 0 0 13 12 0 3
595 575
595 654
705 654
0 1 10 0 0 8192 0 0 13 13 0 3
617 557
617 636
705 636
2 0 11 0 0 8320 0 14 0 0 31 4
704 595
430 595
430 141
500 141
3 1 12 0 0 12416 0 15 14 0 0 4
679 566
686 566
686 577
704 577
0 2 9 0 0 4096 0 0 15 20 0 3
544 449
544 575
630 575
0 1 10 0 0 8320 0 0 15 33 0 5
968 176
968 520
612 520
612 557
630 557
5 3 13 0 0 8320 0 16 25 0 0 4
768 462
857 462
857 194
895 194
3 2 14 0 0 4224 0 17 16 0 0 2
678 458
718 458
0 4 15 0 0 8320 0 0 16 26 0 5
264 368
264 506
711 506
711 476
718 476
1 3 16 0 0 4224 0 6 16 0 0 5
374 84
374 493
693 493
693 467
718 467
0 1 17 0 0 4224 0 0 16 25 0 5
674 322
674 424
698 424
698 449
718 449
0 2 18 0 0 8192 0 0 17 22 0 3
235 396
235 467
633 467
0 1 9 0 0 8192 0 0 17 28 0 3
491 334
491 449
633 449
5 1 19 0 0 8320 0 18 25 0 0 4
749 335
827 335
827 176
895 176
1 4 18 0 0 8320 0 3 18 0 0 5
103 72
103 396
682 396
682 349
699 349
1 3 20 0 0 8320 0 5 18 0 0 5
292 81
292 379
653 379
653 340
699 340
3 2 21 0 0 12416 0 19 18 0 0 4
606 359
635 359
635 331
699 331
3 1 17 0 0 0 0 21 18 0 0 4
649 279
666 279
666 322
699 322
1 2 15 0 0 0 0 4 19 0 0 3
207 73
207 368
561 368
2 1 22 0 0 8320 0 20 19 0 0 4
542 334
554 334
554 350
561 350
0 1 9 0 0 8320 0 0 20 32 0 4
522 167
468 167
468 334
506 334
1 2 5 0 0 0 0 7 21 0 0 3
447 88
447 288
604 288
3 1 23 0 0 4224 0 22 21 0 0 3
593 228
593 270
604 270
1 2 11 0 0 0 0 9 22 0 0 6
576 99
589 99
589 132
500 132
500 237
544 237
1 1 9 0 0 0 0 8 22 0 0 4
511 93
522 93
522 219
544 219
6 1 10 0 0 128 0 25 23 0 0 3
943 176
1114 176
1114 98
1 4 24 0 0 8320 0 2 25 0 0 5
925 286
947 286
947 229
919 229
919 224
10
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1106 29 1143 53
1116 37 1132 53
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
971 25 1024 49
981 33 1013 49
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
852 572 961 596
862 580 950 596
11 Cout and p1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
788 554 841 578
798 562 830 578
4 Cout
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
625 514 702 538
635 522 691 538
7 Q xor B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
728 401 773 425
738 409 762 425
3 KAi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
615 410 660 434
625 418 649 434
3 BP5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
706 276 751 300
716 284 740 300
3 JAi
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
565 302 618 326
575 310 607 326
4 B'P4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
619 221 728 245
629 229 717 245
11 (B xor C)P1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
